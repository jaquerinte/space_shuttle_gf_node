magic
tech gf180mcuC
magscale 1 10
timestamp 1670074230
<< metal1 >>
rect 517346 519374 517358 519426
rect 517410 519423 517422 519426
rect 522498 519423 522510 519426
rect 517410 519377 522510 519423
rect 517410 519374 517422 519377
rect 522498 519374 522510 519377
rect 522562 519374 522574 519426
rect 446898 5966 446910 6018
rect 446962 6015 446974 6018
rect 456194 6015 456206 6018
rect 446962 5969 456206 6015
rect 446962 5966 446974 5969
rect 456194 5966 456206 5969
rect 456258 5966 456270 6018
rect 448802 5854 448814 5906
rect 448866 5903 448878 5906
rect 456306 5903 456318 5906
rect 448866 5857 456318 5903
rect 448866 5854 448878 5857
rect 456306 5854 456318 5857
rect 456370 5854 456382 5906
<< via1 >>
rect 517358 519374 517410 519426
rect 522510 519374 522562 519426
rect 446910 5966 446962 6018
rect 456206 5966 456258 6018
rect 448814 5854 448866 5906
rect 456318 5854 456370 5906
<< metal2 >>
rect 10108 595644 10948 595700
rect 11032 595672 11256 597000
rect 10108 556948 10164 595644
rect 10892 595476 10948 595644
rect 11004 595560 11256 595672
rect 31948 595644 33012 595700
rect 33096 595672 33320 597000
rect 11004 595476 11060 595560
rect 10892 595420 11060 595476
rect 31948 577108 32004 595644
rect 32956 595476 33012 595644
rect 33068 595560 33320 595672
rect 53788 595644 55076 595700
rect 55160 595672 55384 597000
rect 33068 595476 33124 595560
rect 32956 595420 33124 595476
rect 31948 577042 32004 577052
rect 53788 560308 53844 595644
rect 55020 595476 55076 595644
rect 55132 595560 55384 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 99260 595560 99512 595672
rect 121324 595560 121576 595672
rect 142828 595644 143332 595700
rect 143416 595672 143640 597000
rect 55132 595476 55188 595560
rect 55020 595420 55188 595476
rect 53788 560242 53844 560252
rect 10108 556882 10164 556892
rect 5852 556164 5908 556174
rect 2492 547764 2548 547774
rect 140 532644 196 532654
rect 28 521108 84 521118
rect 28 79492 84 521052
rect 140 220612 196 532588
rect 140 220546 196 220556
rect 28 79426 84 79436
rect 2492 51156 2548 547708
rect 2716 534548 2772 534558
rect 2604 527716 2660 527726
rect 2604 305172 2660 527660
rect 2716 403956 2772 534492
rect 5068 524692 5124 524702
rect 5068 516852 5124 524636
rect 5068 516786 5124 516796
rect 2716 403890 2772 403900
rect 2604 305106 2660 305116
rect 5852 107492 5908 556108
rect 17724 554484 17780 554494
rect 12572 547876 12628 547886
rect 9436 542948 9492 542958
rect 9212 542724 9268 542734
rect 5964 537684 6020 537694
rect 5964 192276 6020 537628
rect 6076 519540 6132 519550
rect 6076 262836 6132 519484
rect 6076 262770 6132 262780
rect 5964 192210 6020 192220
rect 5852 107426 5908 107436
rect 9212 93492 9268 542668
rect 9324 529620 9380 529630
rect 9324 418068 9380 529564
rect 9324 418002 9380 418012
rect 9436 333396 9492 542892
rect 10892 541156 10948 541166
rect 9548 521332 9604 521342
rect 9548 502740 9604 521276
rect 9548 502674 9604 502684
rect 9436 333330 9492 333340
rect 10892 248612 10948 541100
rect 11004 537796 11060 537806
rect 11004 276948 11060 537740
rect 11116 531188 11172 531198
rect 11116 389732 11172 531132
rect 11116 389666 11172 389676
rect 11004 276882 11060 276892
rect 10892 248546 10948 248556
rect 12572 121044 12628 547820
rect 15932 546196 15988 546206
rect 14476 539700 14532 539710
rect 14364 532756 14420 532766
rect 12796 527940 12852 527950
rect 12684 526260 12740 526270
rect 12684 346164 12740 526204
rect 12796 445284 12852 527884
rect 12796 445218 12852 445228
rect 14252 522564 14308 522574
rect 12684 346098 12740 346108
rect 12572 120978 12628 120988
rect 9212 93426 9268 93436
rect 14252 63924 14308 522508
rect 14364 176484 14420 532700
rect 14476 361396 14532 539644
rect 14700 536340 14756 536350
rect 14588 522676 14644 522686
rect 14588 473844 14644 522620
rect 14700 487284 14756 536284
rect 14700 487218 14756 487228
rect 14588 473778 14644 473788
rect 14476 361330 14532 361340
rect 14364 176418 14420 176428
rect 15932 134484 15988 546140
rect 17612 531076 17668 531086
rect 16156 526372 16212 526382
rect 16044 524356 16100 524366
rect 16044 290836 16100 524300
rect 16156 431956 16212 526316
rect 16156 431890 16212 431900
rect 16044 290770 16100 290780
rect 17612 205044 17668 531020
rect 17724 233604 17780 554428
rect 70588 552916 70644 552926
rect 26908 552804 26964 552814
rect 19292 549556 19348 549566
rect 17836 538020 17892 538030
rect 17836 317604 17892 537964
rect 17836 317538 17892 317548
rect 17724 233538 17780 233548
rect 17612 204978 17668 204988
rect 19292 149716 19348 549500
rect 19404 544628 19460 544638
rect 19404 163044 19460 544572
rect 19516 527828 19572 527838
rect 19516 374724 19572 527772
rect 26908 519988 26964 552748
rect 40348 551124 40404 551134
rect 35308 546084 35364 546094
rect 35308 537628 35364 546028
rect 35308 537572 35588 537628
rect 32060 529284 32116 529294
rect 32060 519988 32116 529228
rect 26908 519932 27608 519988
rect 31976 519932 32116 519988
rect 35532 519988 35588 537572
rect 40348 519988 40404 551068
rect 53788 544404 53844 544414
rect 53788 537628 53844 544348
rect 53788 537572 53956 537628
rect 44268 536004 44324 536014
rect 44268 519988 44324 535948
rect 50092 524244 50148 524254
rect 50092 519988 50148 524188
rect 53900 519988 53956 537572
rect 66108 530964 66164 530974
rect 58492 525924 58548 525934
rect 58492 519988 58548 525868
rect 63196 520884 63252 520894
rect 63196 519988 63252 520828
rect 35532 519932 36344 519988
rect 40348 519932 40712 519988
rect 44268 519932 45080 519988
rect 49448 519932 50148 519988
rect 53816 519932 53956 519988
rect 58184 519932 58548 519988
rect 62552 519932 63252 519988
rect 66108 519988 66164 530908
rect 70588 519988 70644 552860
rect 77308 550228 77364 595560
rect 99260 572908 99316 595560
rect 121324 572908 121380 595560
rect 99148 572852 99316 572908
rect 120988 572852 121380 572908
rect 99148 570388 99204 572852
rect 99148 570322 99204 570332
rect 77308 550162 77364 550172
rect 84028 551236 84084 551246
rect 75628 549444 75684 549454
rect 75628 537628 75684 549388
rect 75628 537572 75796 537628
rect 75740 519988 75796 537572
rect 66108 519932 66920 519988
rect 70588 519932 71288 519988
rect 75656 519932 75796 519988
rect 79212 534436 79268 534446
rect 79212 519988 79268 534380
rect 84028 519988 84084 551180
rect 119308 541044 119364 541054
rect 109228 539476 109284 539486
rect 97468 539364 97524 539374
rect 97468 537628 97524 539308
rect 109228 537628 109284 539420
rect 119308 537628 119364 540988
rect 97468 537572 97636 537628
rect 109228 537572 109844 537628
rect 119308 537572 119476 537628
rect 88956 520996 89012 521006
rect 88956 519988 89012 520940
rect 97580 519988 97636 537572
rect 106876 526148 106932 526158
rect 106876 519988 106932 526092
rect 79212 519932 80024 519988
rect 84028 519932 84392 519988
rect 88760 519932 89012 519988
rect 97496 519932 97636 519988
rect 106232 519932 106932 519988
rect 109788 519988 109844 537572
rect 115612 527604 115668 527614
rect 115612 519988 115668 527548
rect 119420 519988 119476 537572
rect 120988 523684 121044 572852
rect 142828 546868 142884 595644
rect 143276 595476 143332 595644
rect 143388 595560 143640 595672
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 165480 595560 165732 595672
rect 187544 595560 187796 595672
rect 143388 595476 143444 595560
rect 143276 595420 143444 595476
rect 165676 590212 165732 595560
rect 165676 590146 165732 590156
rect 167132 590212 167188 590222
rect 167132 568708 167188 590156
rect 187740 590212 187796 595560
rect 208348 595644 209524 595700
rect 209608 595672 209832 597000
rect 187740 590146 187796 590156
rect 188972 590212 189028 590222
rect 167132 568642 167188 568652
rect 188972 567028 189028 590156
rect 188972 566962 189028 566972
rect 142828 546802 142884 546812
rect 206668 548548 206724 548558
rect 179788 542836 179844 542846
rect 166348 541268 166404 541278
rect 122668 539588 122724 539598
rect 122668 537628 122724 539532
rect 149548 537908 149604 537918
rect 122668 537572 122948 537628
rect 120988 523618 121044 523628
rect 109788 519932 110600 519988
rect 114968 519932 115668 519988
rect 119336 519932 119476 519988
rect 122892 519988 122948 537572
rect 131628 536228 131684 536238
rect 128716 523572 128772 523582
rect 128716 519988 128772 523516
rect 122892 519932 123704 519988
rect 128072 519932 128772 519988
rect 131628 519988 131684 536172
rect 136108 536116 136164 536126
rect 136108 519988 136164 536060
rect 141260 534660 141316 534670
rect 141260 519988 141316 534604
rect 131628 519932 132440 519988
rect 136108 519932 136808 519988
rect 141176 519932 141316 519988
rect 144732 532868 144788 532878
rect 144732 519988 144788 532812
rect 149548 519988 149604 537852
rect 166348 537628 166404 541212
rect 166348 537572 166628 537628
rect 157948 532980 158004 532990
rect 154476 526036 154532 526046
rect 154476 519988 154532 525980
rect 144732 519932 145544 519988
rect 149548 519932 149912 519988
rect 154280 519932 154532 519988
rect 157948 519988 158004 532924
rect 163660 524580 163716 524590
rect 163660 519988 163716 524524
rect 157948 519932 158648 519988
rect 163016 519932 163716 519988
rect 166572 519988 166628 537572
rect 171388 531300 171444 531310
rect 171388 519988 171444 531244
rect 175308 529508 175364 529518
rect 175308 519988 175364 529452
rect 179788 519988 179844 542780
rect 206668 537628 206724 548492
rect 208348 543508 208404 595644
rect 209468 595476 209524 595644
rect 209580 595560 209832 595672
rect 230188 595644 231588 595700
rect 231672 595672 231896 597000
rect 209580 595476 209636 595560
rect 209468 595420 209636 595476
rect 208348 543442 208404 543452
rect 220892 593124 220948 593134
rect 215068 541828 215124 541838
rect 206668 537572 206836 537628
rect 201628 534324 201684 534334
rect 184940 529732 184996 529742
rect 184940 519988 184996 529676
rect 194236 524468 194292 524478
rect 189756 521220 189812 521230
rect 189756 519988 189812 521164
rect 194236 519988 194292 524412
rect 198156 523348 198212 523358
rect 198156 519988 198212 523292
rect 166572 519932 167384 519988
rect 171388 519932 171752 519988
rect 175308 519932 176120 519988
rect 179788 519932 180488 519988
rect 184856 519932 184996 519988
rect 189224 519932 189812 519988
rect 193592 519932 194292 519988
rect 197960 519932 198212 519988
rect 201628 519988 201684 534268
rect 206780 519988 206836 537572
rect 211596 523460 211652 523470
rect 211596 519988 211652 523404
rect 201628 519932 202328 519988
rect 206696 519932 206836 519988
rect 211064 519932 211652 519988
rect 215068 519988 215124 541772
rect 219884 523236 219940 523246
rect 219884 519988 219940 523180
rect 220892 523236 220948 593068
rect 220892 523170 220948 523180
rect 223468 555268 223524 555278
rect 215068 519932 215432 519988
rect 219800 519932 219940 519988
rect 223468 519988 223524 555212
rect 228508 551908 228564 551918
rect 228508 537628 228564 551852
rect 228508 537572 228676 537628
rect 228620 519988 228676 537572
rect 230188 523796 230244 595644
rect 231532 595476 231588 595644
rect 231644 595560 231896 595672
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 253736 595560 253988 595672
rect 231644 595476 231700 595560
rect 231532 595420 231700 595476
rect 242732 593348 242788 593358
rect 234332 593236 234388 593246
rect 232652 574644 232708 574654
rect 232652 541828 232708 574588
rect 232652 541762 232708 541772
rect 230188 523730 230244 523740
rect 231868 528052 231924 528062
rect 231868 523572 231924 527996
rect 231868 523506 231924 523516
rect 233436 522788 233492 522798
rect 233436 519988 233492 522732
rect 234332 522788 234388 593180
rect 234332 522722 234388 522732
rect 237916 523572 237972 523582
rect 237916 519988 237972 523516
rect 241836 522788 241892 522798
rect 241836 519988 241892 522732
rect 242732 522788 242788 593292
rect 253932 588868 253988 595560
rect 275772 595560 276024 595672
rect 297388 595644 297780 595700
rect 297864 595672 298088 597000
rect 253932 588802 253988 588812
rect 261212 590548 261268 590558
rect 253708 563668 253764 563678
rect 242732 522722 242788 522732
rect 245308 553588 245364 553598
rect 223468 519932 224168 519988
rect 228536 519932 228676 519988
rect 232904 519932 233492 519988
rect 237272 519932 237972 519988
rect 241640 519932 241892 519988
rect 245308 519988 245364 553532
rect 250348 541828 250404 541838
rect 250348 537628 250404 541772
rect 253708 537628 253764 563612
rect 250348 537572 250516 537628
rect 253708 537572 253988 537628
rect 250460 519988 250516 537572
rect 245308 519932 246008 519988
rect 250376 519932 250516 519988
rect 253932 519988 253988 537572
rect 259756 522788 259812 522798
rect 259756 519988 259812 522732
rect 261212 522788 261268 590492
rect 274652 578788 274708 578798
rect 267148 565348 267204 565358
rect 262108 561988 262164 561998
rect 262108 537628 262164 561932
rect 262108 537572 262724 537628
rect 261212 522722 261268 522732
rect 253932 519932 254744 519988
rect 259112 519932 259812 519988
rect 262668 519988 262724 537572
rect 267148 519988 267204 565292
rect 272748 522788 272804 522798
rect 272748 519988 272804 522732
rect 274652 522788 274708 578732
rect 275772 572908 275828 595560
rect 275548 572852 275828 572908
rect 283948 588868 284004 588878
rect 275548 537628 275604 572852
rect 280588 572068 280644 572078
rect 275548 537572 275828 537628
rect 274652 522722 274708 522732
rect 262668 519932 263480 519988
rect 267148 519932 267848 519988
rect 272216 519932 272804 519988
rect 275772 519988 275828 537572
rect 280588 519988 280644 572012
rect 283948 537628 284004 588812
rect 297388 572068 297444 595644
rect 297724 595476 297780 595644
rect 297836 595560 298088 595672
rect 319228 595644 319844 595700
rect 319928 595672 320152 597000
rect 297836 595476 297892 595560
rect 297724 595420 297892 595476
rect 319228 578788 319284 595644
rect 319788 595476 319844 595644
rect 319900 595560 320152 595672
rect 341068 595644 341908 595700
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 319900 595476 319956 595560
rect 319788 595420 319956 595476
rect 319228 578722 319284 578732
rect 335132 590660 335188 590670
rect 297388 572002 297444 572012
rect 332668 577108 332724 577118
rect 319228 570388 319284 570398
rect 305788 568708 305844 568718
rect 297388 567028 297444 567038
rect 288988 543508 289044 543518
rect 283948 537572 284564 537628
rect 284508 519988 284564 537572
rect 288988 519988 289044 543452
rect 297388 537628 297444 566972
rect 302428 546868 302484 546878
rect 297388 537572 297668 537628
rect 294140 523796 294196 523806
rect 294140 519988 294196 523740
rect 275772 519932 276584 519988
rect 280588 519932 280952 519988
rect 284508 519932 285320 519988
rect 288988 519932 289688 519988
rect 294056 519932 294196 519988
rect 297612 519988 297668 537572
rect 302428 519988 302484 546812
rect 305788 537628 305844 568652
rect 315868 550228 315924 550238
rect 315868 537628 315924 550172
rect 319228 537628 319284 570332
rect 324268 560308 324324 560318
rect 305788 537572 306404 537628
rect 315868 537572 316036 537628
rect 319228 537572 319508 537628
rect 306348 519988 306404 537572
rect 310828 523684 310884 523694
rect 310828 519988 310884 523628
rect 315980 519988 316036 537572
rect 297612 519932 298424 519988
rect 302428 519932 302792 519988
rect 306348 519932 307160 519988
rect 310828 519932 311528 519988
rect 315896 519932 316036 519988
rect 319452 519988 319508 537572
rect 324268 519988 324324 560252
rect 327628 556948 327684 556958
rect 327628 537628 327684 556892
rect 327628 537572 328244 537628
rect 328188 519988 328244 537572
rect 332668 519988 332724 577052
rect 335132 565348 335188 590604
rect 335132 565282 335188 565292
rect 337708 586404 337764 586414
rect 337708 537628 337764 586348
rect 341068 561988 341124 595644
rect 341852 595476 341908 595644
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 430220 595560 430472 595672
rect 452284 595560 452536 595672
rect 473788 595644 474292 595700
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 341964 595476 342020 595560
rect 341852 595420 342020 595476
rect 364028 590660 364084 595560
rect 364028 590594 364084 590604
rect 365372 590660 365428 590670
rect 341068 561922 341124 561932
rect 346108 572964 346164 572974
rect 343532 561204 343588 561214
rect 341068 557844 341124 557854
rect 341068 537628 341124 557788
rect 343532 548548 343588 561148
rect 343532 548482 343588 548492
rect 337708 537572 337876 537628
rect 341068 537572 341348 537628
rect 337820 519988 337876 537572
rect 319452 519932 320264 519988
rect 324268 519932 324632 519988
rect 328188 519932 329000 519988
rect 332668 519932 333368 519988
rect 337736 519932 337876 519988
rect 341292 519988 341348 537572
rect 346108 519988 346164 572908
rect 365372 553588 365428 590604
rect 386092 590548 386148 595560
rect 386092 590482 386148 590492
rect 365372 553522 365428 553532
rect 349468 544516 349524 544526
rect 349468 537628 349524 544460
rect 408268 541828 408324 595560
rect 430220 572908 430276 595560
rect 452284 590660 452340 595560
rect 452284 590594 452340 590604
rect 430108 572852 430276 572908
rect 430108 563668 430164 572852
rect 430108 563602 430164 563612
rect 450268 554484 450324 554494
rect 408268 541762 408324 541772
rect 414988 542948 415044 542958
rect 411628 539700 411684 539710
rect 349468 537572 350084 537628
rect 350028 519988 350084 537572
rect 371868 536340 371924 536350
rect 359660 529396 359716 529406
rect 354508 524692 354564 524702
rect 354508 519988 354564 524636
rect 359660 519988 359716 529340
rect 367948 522676 368004 522686
rect 341292 519932 342104 519988
rect 346108 519932 346472 519988
rect 350028 519932 350840 519988
rect 354508 519932 355208 519988
rect 359576 519932 359716 519988
rect 363244 521332 363300 521342
rect 363244 519988 363300 521276
rect 367948 519988 368004 522620
rect 371868 519988 371924 536284
rect 398188 534548 398244 534558
rect 393708 531188 393764 531198
rect 389788 529620 389844 529630
rect 385084 527940 385140 527950
rect 381500 526372 381556 526382
rect 381500 519988 381556 526316
rect 363244 519932 363944 519988
rect 367948 519932 368312 519988
rect 371868 519932 372680 519988
rect 381416 519932 381556 519988
rect 385084 519988 385140 527884
rect 389788 519988 389844 529564
rect 393708 519988 393764 531132
rect 398188 519988 398244 534492
rect 403340 527828 403396 527838
rect 403340 519988 403396 527772
rect 385084 519932 385784 519988
rect 389788 519932 390152 519988
rect 393708 519932 394520 519988
rect 398188 519932 398888 519988
rect 403256 519932 403396 519988
rect 406924 526260 406980 526270
rect 406924 519988 406980 526204
rect 411628 519988 411684 539644
rect 414988 537628 415044 542892
rect 441868 541156 441924 541166
rect 425068 538020 425124 538030
rect 425068 537628 425124 537964
rect 436828 537796 436884 537806
rect 436828 537628 436884 537740
rect 414988 537572 415604 537628
rect 425068 537572 425236 537628
rect 436828 537572 437444 537628
rect 415548 519988 415604 537572
rect 420028 527716 420084 527726
rect 420028 519988 420084 527660
rect 425180 519988 425236 537572
rect 406924 519932 407624 519988
rect 411628 519932 411992 519988
rect 415548 519932 416360 519988
rect 420028 519932 420728 519988
rect 425096 519932 425236 519988
rect 428764 524356 428820 524366
rect 428764 519988 428820 524300
rect 437388 519988 437444 537572
rect 441868 519988 441924 541100
rect 450268 537628 450324 554428
rect 472108 546196 472164 546206
rect 468748 544628 468804 544638
rect 463708 537684 463764 537694
rect 450268 537572 450548 537628
rect 447020 532644 447076 532654
rect 447020 519988 447076 532588
rect 428764 519932 429464 519988
rect 437388 519932 438200 519988
rect 441868 519932 442568 519988
rect 446936 519932 447076 519988
rect 450492 519988 450548 537572
rect 459228 532756 459284 532766
rect 455308 531076 455364 531086
rect 455308 519988 455364 531020
rect 459228 519988 459284 532700
rect 463708 519988 463764 537628
rect 468748 537628 468804 544572
rect 472108 537628 472164 546140
rect 468748 537572 468916 537628
rect 472108 537572 472388 537628
rect 468860 519988 468916 537572
rect 450492 519932 451304 519988
rect 455308 519932 455672 519988
rect 459228 519932 460040 519988
rect 463708 519932 464408 519988
rect 468776 519932 468916 519988
rect 472332 519988 472388 537572
rect 473788 523572 473844 595644
rect 474236 595476 474292 595644
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518476 595560 518728 595672
rect 539308 595644 540484 595700
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 474348 595476 474404 595560
rect 474236 595420 474404 595476
rect 496412 593348 496468 595560
rect 496412 593282 496468 593292
rect 518476 593236 518532 595560
rect 518476 593170 518532 593180
rect 496412 590548 496468 590558
rect 490588 556164 490644 556174
rect 473788 523506 473844 523516
rect 477148 549556 477204 549566
rect 477148 519988 477204 549500
rect 480508 547876 480564 547886
rect 480508 537628 480564 547820
rect 485548 542724 485604 542734
rect 480508 537572 481124 537628
rect 481068 519988 481124 537572
rect 485548 519988 485604 542668
rect 490588 537628 490644 556108
rect 496412 551908 496468 590492
rect 539308 555268 539364 595644
rect 540428 595476 540484 595644
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 540540 595476 540596 595560
rect 540428 595420 540596 595476
rect 562604 590548 562660 595560
rect 584668 593124 584724 595560
rect 584668 593058 584724 593068
rect 562604 590482 562660 590492
rect 539308 555202 539364 555212
rect 590604 588644 590660 588654
rect 496412 551842 496468 551852
rect 568652 552916 568708 552926
rect 498988 547764 499044 547774
rect 490588 537572 490756 537628
rect 490700 519988 490756 537572
rect 472332 519932 473144 519988
rect 477148 519932 477512 519988
rect 481068 519932 481880 519988
rect 485548 519932 486248 519988
rect 490616 519932 490756 519988
rect 494284 521108 494340 521118
rect 494284 519988 494340 521052
rect 498988 519988 499044 547708
rect 526652 544404 526708 544414
rect 521612 534660 521668 534670
rect 513100 522788 513156 522798
rect 508732 522676 508788 522686
rect 503020 522564 503076 522574
rect 503020 519988 503076 522508
rect 508732 519988 508788 522620
rect 513100 519988 513156 522732
rect 494284 519932 494984 519988
rect 498988 519932 499352 519988
rect 503020 519932 503720 519988
rect 508088 519932 508788 519988
rect 512456 519932 513156 519988
rect 519372 522676 519428 522686
rect 19628 519652 19684 519662
rect 19628 458724 19684 519596
rect 377020 519652 377076 519662
rect 377020 519586 377076 519596
rect 433804 519540 433860 519550
rect 433804 519474 433860 519484
rect 93100 519428 93156 519438
rect 517356 519428 517412 519438
rect 516824 519426 517412 519428
rect 516824 519374 517358 519426
rect 517410 519374 517412 519426
rect 516824 519372 517412 519374
rect 93100 519362 93156 519372
rect 517356 519362 517412 519372
rect 23212 519316 23268 519326
rect 23212 519250 23268 519260
rect 101836 519316 101892 519326
rect 101836 519250 101892 519260
rect 19628 458658 19684 458668
rect 19516 374658 19572 374668
rect 19404 162978 19460 162988
rect 19292 149650 19348 149660
rect 15932 134418 15988 134428
rect 14252 63858 14308 63868
rect 2492 51090 2548 51100
rect 4172 36820 4228 36830
rect 4172 20020 4228 36764
rect 4956 22708 5012 22718
rect 4956 20132 5012 22652
rect 4956 20066 5012 20076
rect 33740 20076 34720 20132
rect 35644 20076 36288 20132
rect 37212 20076 37856 20132
rect 38780 20076 39424 20132
rect 40348 20076 40992 20132
rect 42028 20076 42560 20132
rect 43932 20076 44128 20132
rect 45388 20076 45696 20132
rect 47068 20076 47264 20132
rect 48748 20076 48832 20132
rect 4172 19954 4228 19964
rect 32732 18340 32788 18350
rect 18508 17668 18564 17678
rect 15148 12628 15204 12638
rect 13356 10948 13412 10958
rect 11564 7588 11620 7598
rect 11564 480 11620 7532
rect 13356 480 13412 10892
rect 15148 480 15204 12572
rect 17276 4228 17332 4238
rect 17276 480 17332 4172
rect 11368 392 11620 480
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15148 392 15400 480
rect 15176 -960 15400 392
rect 17080 392 17332 480
rect 18508 420 18564 17612
rect 30380 15988 30436 15998
rect 22988 5908 23044 5918
rect 21084 4340 21140 4350
rect 18844 480 19012 532
rect 21084 480 21140 4284
rect 22988 480 23044 5852
rect 28700 4676 28756 4686
rect 24892 4564 24948 4574
rect 24892 480 24948 4508
rect 26796 4452 26852 4462
rect 26796 480 26852 4396
rect 28700 480 28756 4620
rect 18844 476 19208 480
rect 18844 420 18900 476
rect 17080 -960 17304 392
rect 18508 364 18900 420
rect 18956 392 19208 476
rect 18984 -960 19208 392
rect 20888 392 21140 480
rect 22792 392 23044 480
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 28504 392 28756 480
rect 30380 480 30436 15932
rect 31948 14308 32004 14318
rect 30380 392 30632 480
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 31948 420 32004 14252
rect 32732 5908 32788 18284
rect 32732 5842 32788 5852
rect 33628 18116 33684 18126
rect 32172 480 32340 532
rect 32172 476 32536 480
rect 32172 420 32228 476
rect 31948 364 32228 420
rect 32284 392 32536 476
rect 32312 -960 32536 392
rect 33628 420 33684 18060
rect 33740 7588 33796 20076
rect 33740 7522 33796 7532
rect 35308 18004 35364 18014
rect 34076 480 34244 532
rect 34076 476 34440 480
rect 34076 420 34132 476
rect 33628 364 34132 420
rect 34188 392 34440 476
rect 34216 -960 34440 392
rect 35308 420 35364 17948
rect 35644 10948 35700 20076
rect 35644 10882 35700 10892
rect 36988 17892 37044 17902
rect 35980 480 36148 532
rect 35980 476 36344 480
rect 35980 420 36036 476
rect 35308 364 36036 420
rect 36092 392 36344 476
rect 36120 -960 36344 392
rect 36988 420 37044 17836
rect 37212 12628 37268 20076
rect 37212 12562 37268 12572
rect 38668 17780 38724 17790
rect 37884 480 38052 532
rect 37884 476 38248 480
rect 37884 420 37940 476
rect 36988 364 37940 420
rect 37996 392 38248 476
rect 38024 -960 38248 392
rect 38668 420 38724 17724
rect 38780 4228 38836 20076
rect 40348 17668 40404 20076
rect 40348 17602 40404 17612
rect 40460 18228 40516 18238
rect 38780 4162 38836 4172
rect 39788 480 39956 532
rect 39788 476 40152 480
rect 39788 420 39844 476
rect 38668 364 39844 420
rect 39900 392 40152 476
rect 39928 -960 40152 392
rect 40460 420 40516 18172
rect 42028 4340 42084 20076
rect 43932 18340 43988 20076
rect 43932 18274 43988 18284
rect 42028 4274 42084 4284
rect 43932 11060 43988 11070
rect 41692 480 41860 532
rect 43932 480 43988 11004
rect 45388 4564 45444 20076
rect 45388 4498 45444 4508
rect 45836 11620 45892 11630
rect 45836 480 45892 11564
rect 47068 4452 47124 20076
rect 47068 4386 47124 4396
rect 47740 11284 47796 11294
rect 47740 480 47796 11228
rect 48748 4676 48804 20076
rect 50428 15988 50484 20104
rect 50428 15922 50484 15932
rect 51324 20076 51968 20132
rect 52892 20076 53536 20132
rect 54460 20076 55104 20132
rect 56364 20076 56672 20132
rect 57596 20076 58240 20132
rect 59164 20076 59808 20132
rect 60732 20076 61376 20132
rect 62300 20076 62944 20132
rect 63980 20076 64512 20132
rect 65660 20076 66080 20132
rect 67452 20076 67648 20132
rect 68908 20076 69216 20132
rect 70588 20076 70784 20132
rect 72268 20076 72352 20132
rect 73976 20076 74340 20132
rect 51324 14308 51380 20076
rect 52892 18116 52948 20076
rect 52892 18050 52948 18060
rect 54460 18004 54516 20076
rect 54460 17938 54516 17948
rect 56364 17892 56420 20076
rect 56364 17826 56420 17836
rect 57596 17780 57652 20076
rect 59164 18228 59220 20076
rect 59164 18162 59220 18172
rect 57596 17714 57652 17724
rect 51324 14242 51380 14252
rect 60508 17668 60564 17678
rect 48748 4610 48804 4620
rect 49644 11508 49700 11518
rect 49644 480 49700 11452
rect 55356 11396 55412 11406
rect 51548 11172 51604 11182
rect 51548 480 51604 11116
rect 53452 10948 53508 10958
rect 53452 480 53508 10892
rect 55356 480 55412 11340
rect 57260 4340 57316 4350
rect 57260 480 57316 4284
rect 59164 4228 59220 4238
rect 59164 480 59220 4172
rect 41692 476 42056 480
rect 41692 420 41748 476
rect 40460 364 41748 420
rect 41804 392 42056 476
rect 41832 -960 42056 392
rect 43736 392 43988 480
rect 45640 392 45892 480
rect 47544 392 47796 480
rect 49448 392 49700 480
rect 51352 392 51604 480
rect 53256 392 53508 480
rect 55160 392 55412 480
rect 57064 392 57316 480
rect 58968 392 59220 480
rect 60508 420 60564 17612
rect 60732 11060 60788 20076
rect 60732 10994 60788 11004
rect 62188 17892 62244 17902
rect 60732 480 60900 532
rect 60732 476 61096 480
rect 60732 420 60788 476
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 392
rect 53256 -960 53480 392
rect 55160 -960 55384 392
rect 57064 -960 57288 392
rect 58968 -960 59192 392
rect 60508 364 60788 420
rect 60844 392 61096 476
rect 60872 -960 61096 392
rect 62188 420 62244 17836
rect 62300 11620 62356 20076
rect 62300 11554 62356 11564
rect 63868 18004 63924 18014
rect 62636 480 62804 532
rect 62636 476 63000 480
rect 62636 420 62692 476
rect 62188 364 62692 420
rect 62748 392 63000 476
rect 62776 -960 63000 392
rect 63868 420 63924 17948
rect 63980 11284 64036 20076
rect 63980 11218 64036 11228
rect 65548 17780 65604 17790
rect 64540 480 64708 532
rect 64540 476 64904 480
rect 64540 420 64596 476
rect 63868 364 64596 420
rect 64652 392 64904 476
rect 64680 -960 64904 392
rect 65548 420 65604 17724
rect 65660 11508 65716 20076
rect 65660 11442 65716 11452
rect 67228 18116 67284 18126
rect 66444 480 66612 532
rect 66444 476 66808 480
rect 66444 420 66500 476
rect 65548 364 66500 420
rect 66556 392 66808 476
rect 66584 -960 66808 392
rect 67228 420 67284 18060
rect 67452 11172 67508 20076
rect 67452 11106 67508 11116
rect 68908 10948 68964 20076
rect 68908 10882 68964 10892
rect 69020 18228 69076 18238
rect 69020 8428 69076 18172
rect 70588 11396 70644 20076
rect 70588 11330 70644 11340
rect 68908 8372 69076 8428
rect 68348 480 68516 532
rect 68348 476 68712 480
rect 68348 420 68404 476
rect 67228 364 68404 420
rect 68460 392 68712 476
rect 68488 -960 68712 392
rect 68908 420 68964 8372
rect 72268 4340 72324 20076
rect 72268 4274 72324 4284
rect 72380 13300 72436 13310
rect 70252 480 70420 532
rect 72380 480 72436 13244
rect 74172 13188 74228 13198
rect 74172 480 74228 13132
rect 74284 4228 74340 20076
rect 74844 20076 75488 20132
rect 76412 20076 77056 20132
rect 77980 20076 78624 20132
rect 79884 20076 80192 20132
rect 81116 20076 81760 20132
rect 82684 20076 83328 20132
rect 84252 20076 84896 20132
rect 85820 20076 86464 20132
rect 87388 20076 88032 20132
rect 89180 20076 89600 20132
rect 90972 20076 91168 20132
rect 92428 20076 92736 20132
rect 94220 20076 94304 20132
rect 95788 20076 95872 20132
rect 74844 17668 74900 20076
rect 76412 17892 76468 20076
rect 77980 18004 78036 20076
rect 77980 17938 78036 17948
rect 76412 17826 76468 17836
rect 79884 17780 79940 20076
rect 81116 18116 81172 20076
rect 82684 18228 82740 20076
rect 82684 18162 82740 18172
rect 81116 18050 81172 18060
rect 79884 17714 79940 17724
rect 74844 17602 74900 17612
rect 84252 13300 84308 20076
rect 84252 13234 84308 13244
rect 85708 17780 85764 17790
rect 80668 13076 80724 13086
rect 77308 12852 77364 12862
rect 74284 4162 74340 4172
rect 75628 12740 75684 12750
rect 70252 476 70616 480
rect 70252 420 70308 476
rect 68908 364 70308 420
rect 70364 392 70616 476
rect 70392 -960 70616 392
rect 72296 -960 72520 480
rect 74172 392 74424 480
rect 74200 -960 74424 392
rect 75628 420 75684 12684
rect 75964 480 76132 532
rect 75964 476 76328 480
rect 75964 420 76020 476
rect 75628 364 76020 420
rect 76076 392 76328 476
rect 76104 -960 76328 392
rect 77308 420 77364 12796
rect 78988 12628 79044 12638
rect 77868 480 78036 532
rect 77868 476 78232 480
rect 77868 420 77924 476
rect 77308 364 77924 420
rect 77980 392 78232 476
rect 78008 -960 78232 392
rect 78988 420 79044 12572
rect 79772 480 79940 532
rect 79772 476 80136 480
rect 79772 420 79828 476
rect 78988 364 79828 420
rect 79884 392 80136 476
rect 79912 -960 80136 392
rect 80668 420 80724 13020
rect 82348 12964 82404 12974
rect 81676 480 81844 532
rect 81676 476 82040 480
rect 81676 420 81732 476
rect 80668 364 81732 420
rect 81788 392 82040 476
rect 81816 -960 82040 392
rect 82348 420 82404 12908
rect 83580 480 83748 532
rect 85708 480 85764 17724
rect 85820 13188 85876 20076
rect 85820 13122 85876 13132
rect 87388 12740 87444 20076
rect 89068 18004 89124 18014
rect 87388 12674 87444 12684
rect 87500 17668 87556 17678
rect 87500 480 87556 17612
rect 83580 476 83944 480
rect 83580 420 83636 476
rect 82348 364 83636 420
rect 83692 392 83944 476
rect 83720 -960 83944 392
rect 85624 -960 85848 480
rect 87500 392 87752 480
rect 87528 -960 87752 392
rect 89068 420 89124 17948
rect 89180 12852 89236 20076
rect 89180 12786 89236 12796
rect 90748 18228 90804 18238
rect 89292 480 89460 532
rect 89292 476 89656 480
rect 89292 420 89348 476
rect 89068 364 89348 420
rect 89404 392 89656 476
rect 89432 -960 89656 392
rect 90748 420 90804 18172
rect 90972 12628 91028 20076
rect 92428 13076 92484 20076
rect 92428 13010 92484 13020
rect 92540 18340 92596 18350
rect 90972 12562 91028 12572
rect 92540 8428 92596 18284
rect 92428 8372 92596 8428
rect 94108 16996 94164 17006
rect 91196 480 91364 532
rect 91196 476 91560 480
rect 91196 420 91252 476
rect 90748 364 91252 420
rect 91308 392 91560 476
rect 91336 -960 91560 392
rect 92428 420 92484 8372
rect 93100 480 93268 532
rect 93100 476 93464 480
rect 93100 420 93156 476
rect 92428 364 93156 420
rect 93212 392 93464 476
rect 93240 -960 93464 392
rect 94108 420 94164 16940
rect 94220 12964 94276 20076
rect 95788 17780 95844 20076
rect 95788 17714 95844 17724
rect 97468 17668 97524 20104
rect 98364 20076 99008 20132
rect 99932 20076 100576 20132
rect 101500 20076 102144 20132
rect 103516 20076 103712 20132
rect 104636 20076 105280 20132
rect 106204 20076 106848 20132
rect 107772 20076 108416 20132
rect 109340 20076 109984 20132
rect 110908 20076 111552 20132
rect 112588 20076 113120 20132
rect 114492 20076 114688 20132
rect 115948 20076 116256 20132
rect 117628 20076 117824 20132
rect 119308 20076 119392 20132
rect 97468 17602 97524 17612
rect 97692 18452 97748 18462
rect 94220 12898 94276 12908
rect 95900 16884 95956 16894
rect 95004 480 95172 532
rect 95004 476 95368 480
rect 95004 420 95060 476
rect 94108 364 95060 420
rect 95116 392 95368 476
rect 95144 -960 95368 392
rect 95900 420 95956 16828
rect 96908 480 97076 532
rect 96908 476 97272 480
rect 96908 420 96964 476
rect 95900 364 96964 420
rect 97020 392 97272 476
rect 97048 -960 97272 392
rect 97692 420 97748 18396
rect 98364 18004 98420 20076
rect 99932 18228 99988 20076
rect 101500 18340 101556 20076
rect 101500 18274 101556 18284
rect 99932 18162 99988 18172
rect 98364 17938 98420 17948
rect 102732 18116 102788 18126
rect 100828 17668 100884 17678
rect 98812 480 98980 532
rect 100828 480 100884 17612
rect 102732 480 102788 18060
rect 103516 16996 103572 20076
rect 103516 16930 103572 16940
rect 104188 18004 104244 18014
rect 98812 476 99176 480
rect 98812 420 98868 476
rect 97692 364 98868 420
rect 98924 392 99176 476
rect 100828 392 101080 480
rect 102732 392 102984 480
rect 98952 -960 99176 392
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104188 420 104244 17948
rect 104636 16884 104692 20076
rect 106204 18452 106260 20076
rect 106204 18386 106260 18396
rect 104636 16818 104692 16828
rect 105868 18228 105924 18238
rect 104524 480 104692 532
rect 104524 476 104888 480
rect 104524 420 104580 476
rect 104188 364 104580 420
rect 104636 392 104888 476
rect 104664 -960 104888 392
rect 105868 420 105924 18172
rect 107772 17668 107828 20076
rect 109340 18116 109396 20076
rect 109340 18050 109396 18060
rect 110908 18004 110964 20076
rect 112588 18228 112644 20076
rect 112588 18162 112644 18172
rect 110908 17938 110964 17948
rect 107772 17602 107828 17612
rect 110908 17780 110964 17790
rect 107660 16996 107716 17006
rect 106428 480 106596 532
rect 106428 476 106792 480
rect 106428 420 106484 476
rect 105868 364 106484 420
rect 106540 392 106792 476
rect 106568 -960 106792 392
rect 107660 420 107716 16940
rect 109228 16884 109284 16894
rect 108332 480 108500 532
rect 108332 476 108696 480
rect 108332 420 108388 476
rect 107660 364 108388 420
rect 108444 392 108696 476
rect 108472 -960 108696 392
rect 109228 420 109284 16828
rect 110236 480 110404 532
rect 110236 476 110600 480
rect 110236 420 110292 476
rect 109228 364 110292 420
rect 110348 392 110600 476
rect 110376 -960 110600 392
rect 110908 420 110964 17724
rect 114268 17668 114324 17678
rect 112140 480 112308 532
rect 114268 480 114324 17612
rect 114492 16996 114548 20076
rect 114492 16930 114548 16940
rect 115948 16884 116004 20076
rect 117628 17780 117684 20076
rect 117628 17714 117684 17724
rect 119308 17668 119364 20076
rect 119308 17602 119364 17612
rect 115948 16818 116004 16828
rect 116060 16996 116116 17006
rect 116060 480 116116 16940
rect 120988 16996 121044 20104
rect 120988 16930 121044 16940
rect 121884 20076 122528 20132
rect 123452 20076 124096 20132
rect 125020 20076 125664 20132
rect 126924 20076 127232 20132
rect 128156 20076 128800 20132
rect 129724 20076 130368 20132
rect 131404 20076 131936 20132
rect 132860 20076 133504 20132
rect 134428 20076 135072 20132
rect 136108 20076 136640 20132
rect 138012 20076 138208 20132
rect 139580 20076 139776 20132
rect 141148 20076 141344 20132
rect 142828 20076 142912 20132
rect 144536 20076 144676 20132
rect 117628 15092 117684 15102
rect 112140 476 112504 480
rect 112140 420 112196 476
rect 110908 364 112196 420
rect 112252 392 112504 476
rect 112280 -960 112504 392
rect 114184 -960 114408 480
rect 116060 392 116312 480
rect 116088 -960 116312 392
rect 117628 420 117684 15036
rect 121884 15092 121940 20076
rect 121884 15026 121940 15036
rect 122780 15092 122836 15102
rect 120988 14980 121044 14990
rect 119308 14756 119364 14766
rect 117852 480 118020 532
rect 117852 476 118216 480
rect 117852 420 117908 476
rect 117628 364 117908 420
rect 117964 392 118216 476
rect 117992 -960 118216 392
rect 119308 420 119364 14700
rect 119756 480 119924 532
rect 119756 476 120120 480
rect 119756 420 119812 476
rect 119308 364 119812 420
rect 119868 392 120120 476
rect 119896 -960 120120 392
rect 120988 420 121044 14924
rect 121660 480 121828 532
rect 121660 476 122024 480
rect 121660 420 121716 476
rect 120988 364 121716 420
rect 121772 392 122024 476
rect 121800 -960 122024 392
rect 122780 420 122836 15036
rect 123452 14756 123508 20076
rect 125020 14980 125076 20076
rect 126924 15092 126980 20076
rect 126924 15026 126980 15036
rect 125020 14914 125076 14924
rect 123452 14690 123508 14700
rect 126028 14868 126084 14878
rect 124348 14420 124404 14430
rect 123564 480 123732 532
rect 123564 476 123928 480
rect 123564 420 123620 476
rect 122780 364 123620 420
rect 123676 392 123928 476
rect 123704 -960 123928 392
rect 124348 420 124404 14364
rect 125468 480 125636 532
rect 125468 476 125832 480
rect 125468 420 125524 476
rect 124348 364 125524 420
rect 125580 392 125832 476
rect 125608 -960 125832 392
rect 126028 420 126084 14812
rect 128156 14420 128212 20076
rect 129724 14868 129780 20076
rect 129724 14802 129780 14812
rect 128156 14354 128212 14364
rect 131292 13412 131348 13422
rect 129388 13300 129444 13310
rect 127372 480 127540 532
rect 129388 480 129444 13244
rect 131292 480 131348 13356
rect 131404 13300 131460 20076
rect 132860 13412 132916 20076
rect 132860 13346 132916 13356
rect 131404 13234 131460 13244
rect 132748 13300 132804 13310
rect 127372 476 127736 480
rect 127372 420 127428 476
rect 126028 364 127428 420
rect 127484 392 127736 476
rect 129388 392 129640 480
rect 131292 392 131544 480
rect 127512 -960 127736 392
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 132748 420 132804 13244
rect 134428 13300 134484 20076
rect 134428 13234 134484 13244
rect 134540 13412 134596 13422
rect 133084 480 133252 532
rect 133084 476 133448 480
rect 133084 420 133140 476
rect 132748 364 133140 420
rect 133196 392 133448 476
rect 133224 -960 133448 392
rect 134540 420 134596 13356
rect 136108 13412 136164 20076
rect 136108 13346 136164 13356
rect 137900 13300 137956 13310
rect 136108 12068 136164 12078
rect 134988 480 135156 532
rect 134988 476 135352 480
rect 134988 420 135044 476
rect 134540 364 135044 420
rect 135100 392 135352 476
rect 135128 -960 135352 392
rect 136108 420 136164 12012
rect 136892 480 137060 532
rect 136892 476 137256 480
rect 136892 420 136948 476
rect 136108 364 136948 420
rect 137004 392 137256 476
rect 137032 -960 137256 392
rect 137900 420 137956 13244
rect 138012 12068 138068 20076
rect 138012 12002 138068 12012
rect 139468 13412 139524 13422
rect 138796 480 138964 532
rect 138796 476 139160 480
rect 138796 420 138852 476
rect 137900 364 138852 420
rect 138908 392 139160 476
rect 138936 -960 139160 392
rect 139468 420 139524 13356
rect 139580 13300 139636 20076
rect 141148 13412 141204 20076
rect 141148 13346 141204 13356
rect 139580 13234 139636 13244
rect 140700 480 140868 532
rect 142828 480 142884 20076
rect 144620 480 144676 20076
rect 144732 20076 146048 20132
rect 146188 20076 147616 20132
rect 147868 20076 149184 20132
rect 149548 20076 150752 20132
rect 151228 20076 152320 20132
rect 152908 20076 153888 20132
rect 154588 20076 155456 20132
rect 156268 20076 157024 20132
rect 158060 20076 158592 20132
rect 159628 20076 160160 20132
rect 161308 20076 161728 20132
rect 162988 20076 163296 20132
rect 164668 20076 164864 20132
rect 166348 20076 166432 20132
rect 144732 4676 144788 20076
rect 144732 4610 144788 4620
rect 146188 4340 146244 20076
rect 147868 5012 147924 20076
rect 147868 4946 147924 4956
rect 146188 4274 146244 4284
rect 146524 4676 146580 4686
rect 146524 480 146580 4620
rect 148428 4340 148484 4350
rect 148428 480 148484 4284
rect 149548 4340 149604 20076
rect 149548 4274 149604 4284
rect 150332 5012 150388 5022
rect 150332 480 150388 4956
rect 151228 4228 151284 20076
rect 151228 4162 151284 4172
rect 152236 4340 152292 4350
rect 152236 480 152292 4284
rect 152908 4340 152964 20076
rect 154588 4676 154644 20076
rect 154588 4610 154644 4620
rect 152908 4274 152964 4284
rect 156044 4340 156100 4350
rect 154140 4228 154196 4238
rect 154140 480 154196 4172
rect 156044 480 156100 4284
rect 156268 4228 156324 20076
rect 158060 4788 158116 20076
rect 159628 4900 159684 20076
rect 159628 4834 159684 4844
rect 158060 4722 158116 4732
rect 156268 4162 156324 4172
rect 157948 4676 158004 4686
rect 157948 480 158004 4620
rect 159852 4228 159908 4238
rect 159852 480 159908 4172
rect 161308 4228 161364 20076
rect 161308 4162 161364 4172
rect 161756 4788 161812 4798
rect 161756 480 161812 4732
rect 162988 4340 163044 20076
rect 162988 4274 163044 4284
rect 163660 4900 163716 4910
rect 163660 480 163716 4844
rect 164668 4116 164724 20076
rect 166348 4564 166404 20076
rect 168028 4788 168084 20104
rect 168140 20076 169568 20132
rect 169708 20076 171136 20132
rect 171388 20076 172704 20132
rect 173068 20076 174272 20132
rect 174748 20076 175840 20132
rect 176428 20076 177408 20132
rect 178108 20076 178976 20132
rect 179788 20076 180544 20132
rect 181468 20076 182112 20132
rect 183148 20076 183680 20132
rect 184828 20076 185248 20132
rect 186508 20076 186816 20132
rect 188188 20076 188384 20132
rect 189868 20076 189952 20132
rect 168140 6020 168196 20076
rect 168140 5954 168196 5964
rect 169708 5908 169764 20076
rect 171388 6132 171444 20076
rect 171388 6066 171444 6076
rect 169708 5842 169764 5852
rect 173068 5124 173124 20076
rect 174748 6244 174804 20076
rect 176428 6468 176484 20076
rect 176428 6402 176484 6412
rect 174748 6178 174804 6188
rect 173068 5058 173124 5068
rect 175084 6020 175140 6030
rect 168028 4722 168084 4732
rect 173180 4788 173236 4798
rect 166348 4498 166404 4508
rect 171388 4564 171444 4574
rect 167468 4340 167524 4350
rect 164668 4050 164724 4060
rect 165564 4228 165620 4238
rect 165564 480 165620 4172
rect 167468 480 167524 4284
rect 169372 4116 169428 4126
rect 169372 480 169428 4060
rect 171388 480 171444 4508
rect 173180 480 173236 4732
rect 175084 480 175140 5964
rect 176988 5908 177044 5918
rect 176988 480 177044 5852
rect 178108 5796 178164 20076
rect 178108 5730 178164 5740
rect 178892 6132 178948 6142
rect 178892 480 178948 6076
rect 179788 5908 179844 20076
rect 181468 6132 181524 20076
rect 181468 6066 181524 6076
rect 182700 6244 182756 6254
rect 179788 5842 179844 5852
rect 180796 5124 180852 5134
rect 180796 480 180852 5068
rect 182700 480 182756 6188
rect 183148 6244 183204 20076
rect 183148 6178 183204 6188
rect 184604 6468 184660 6478
rect 184604 480 184660 6412
rect 184828 5124 184884 20076
rect 186508 6356 186564 20076
rect 186508 6290 186564 6300
rect 188188 6020 188244 20076
rect 188188 5954 188244 5964
rect 188412 5908 188468 5918
rect 184828 5058 184884 5068
rect 186508 5796 186564 5806
rect 186508 480 186564 5740
rect 188412 480 188468 5852
rect 189868 4228 189924 20076
rect 189868 4162 189924 4172
rect 190316 6132 190372 6142
rect 190316 480 190372 6076
rect 191548 4340 191604 20104
rect 191660 20076 193088 20132
rect 193228 20076 194656 20132
rect 194908 20076 196224 20132
rect 196588 20076 197792 20132
rect 198268 20076 199360 20132
rect 199948 20076 200928 20132
rect 191660 6468 191716 20076
rect 191660 6402 191716 6412
rect 191548 4274 191604 4284
rect 192220 6244 192276 6254
rect 192220 480 192276 6188
rect 193228 6020 193284 20076
rect 194908 6244 194964 20076
rect 194908 6178 194964 6188
rect 196028 6356 196084 6366
rect 193228 5954 193284 5964
rect 194124 5124 194180 5134
rect 194124 480 194180 5068
rect 196028 480 196084 6300
rect 196588 6356 196644 20076
rect 196588 6290 196644 6300
rect 198268 6132 198324 20076
rect 198268 6066 198324 6076
rect 197932 5908 197988 5918
rect 197932 480 197988 5852
rect 199948 5908 200004 20076
rect 202524 10948 202580 20104
rect 204092 11284 204148 20104
rect 204092 11218 204148 11228
rect 205660 11060 205716 20104
rect 207228 11620 207284 20104
rect 207228 11554 207284 11564
rect 208796 11172 208852 20104
rect 210364 11396 210420 20104
rect 211932 11508 211988 20104
rect 211932 11442 211988 11452
rect 213388 20076 213472 20132
rect 215096 20076 215236 20132
rect 210364 11330 210420 11340
rect 208796 11106 208852 11116
rect 205660 10994 205716 11004
rect 202524 10882 202580 10892
rect 199948 5842 200004 5852
rect 203644 6468 203700 6478
rect 201740 4340 201796 4350
rect 199948 4228 200004 4238
rect 199948 480 200004 4172
rect 201740 480 201796 4284
rect 203644 480 203700 6412
rect 209356 6356 209412 6366
rect 207452 6244 207508 6254
rect 205548 6020 205604 6030
rect 205548 480 205604 5964
rect 207452 480 207508 6188
rect 209356 480 209412 6300
rect 211260 6132 211316 6142
rect 211260 480 211316 6076
rect 213164 5908 213220 5918
rect 213164 480 213220 5852
rect 213388 5908 213444 20076
rect 213388 5842 213444 5852
rect 215068 10948 215124 10958
rect 215068 480 215124 10892
rect 215180 6020 215236 20076
rect 216636 16548 216692 20104
rect 216636 16482 216692 16492
rect 218204 16100 218260 20104
rect 218204 16034 218260 16044
rect 219772 15988 219828 20104
rect 221340 16324 221396 20104
rect 221340 16258 221396 16268
rect 222908 16212 222964 20104
rect 224476 16436 224532 20104
rect 224476 16370 224532 16380
rect 222908 16146 222964 16156
rect 219772 15922 219828 15932
rect 226044 14308 226100 20104
rect 227612 14532 227668 20104
rect 229180 14644 229236 20104
rect 229180 14578 229236 14588
rect 227612 14466 227668 14476
rect 230748 14420 230804 20104
rect 230748 14354 230804 14364
rect 231868 16548 231924 16558
rect 226044 14242 226100 14252
rect 220780 11620 220836 11630
rect 215180 5954 215236 5964
rect 216972 11284 217028 11294
rect 216972 480 217028 11228
rect 218876 11060 218932 11070
rect 218876 480 218932 11004
rect 220780 480 220836 11564
rect 226492 11508 226548 11518
rect 224588 11396 224644 11406
rect 222684 11172 222740 11182
rect 222684 480 222740 11116
rect 224588 480 224644 11340
rect 226492 480 226548 11452
rect 230300 6020 230356 6030
rect 228508 5908 228564 5918
rect 228508 480 228564 5852
rect 230300 480 230356 5964
rect 140700 476 141064 480
rect 140700 420 140756 476
rect 139468 364 140756 420
rect 140812 392 141064 476
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144620 392 144872 480
rect 146524 392 146776 480
rect 148428 392 148680 480
rect 150332 392 150584 480
rect 152236 392 152488 480
rect 154140 392 154392 480
rect 156044 392 156296 480
rect 157948 392 158200 480
rect 159852 392 160104 480
rect 161756 392 162008 480
rect 163660 392 163912 480
rect 165564 392 165816 480
rect 167468 392 167720 480
rect 169372 392 169624 480
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 392
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173180 392 173432 480
rect 175084 392 175336 480
rect 176988 392 177240 480
rect 178892 392 179144 480
rect 180796 392 181048 480
rect 182700 392 182952 480
rect 184604 392 184856 480
rect 186508 392 186760 480
rect 188412 392 188664 480
rect 190316 392 190568 480
rect 192220 392 192472 480
rect 194124 392 194376 480
rect 196028 392 196280 480
rect 197932 392 198184 480
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 392
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 203644 392 203896 480
rect 205548 392 205800 480
rect 207452 392 207704 480
rect 209356 392 209608 480
rect 211260 392 211512 480
rect 213164 392 213416 480
rect 215068 392 215320 480
rect 216972 392 217224 480
rect 218876 392 219128 480
rect 220780 392 221032 480
rect 222684 392 222936 480
rect 224588 392 224840 480
rect 226492 392 226744 480
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 392
rect 215096 -960 215320 392
rect 217000 -960 217224 392
rect 218904 -960 219128 392
rect 220808 -960 221032 392
rect 222712 -960 222936 392
rect 224616 -960 224840 392
rect 226520 -960 226744 392
rect 228424 -960 228648 480
rect 230300 392 230552 480
rect 230328 -960 230552 392
rect 231868 420 231924 16492
rect 232316 14756 232372 20104
rect 232316 14690 232372 14700
rect 233548 16100 233604 16110
rect 232092 480 232260 532
rect 232092 476 232456 480
rect 232092 420 232148 476
rect 231868 364 232148 420
rect 232204 392 232456 476
rect 232232 -960 232456 392
rect 233548 420 233604 16044
rect 233884 14868 233940 20104
rect 233884 14802 233940 14812
rect 235228 15988 235284 15998
rect 233996 480 234164 532
rect 233996 476 234360 480
rect 233996 420 234052 476
rect 233548 364 234052 420
rect 234108 392 234360 476
rect 234136 -960 234360 392
rect 235228 420 235284 15932
rect 235452 14980 235508 20104
rect 235452 14914 235508 14924
rect 236908 16324 236964 16334
rect 235900 480 236068 532
rect 235900 476 236264 480
rect 235900 420 235956 476
rect 235228 364 235956 420
rect 236012 392 236264 476
rect 236040 -960 236264 392
rect 236908 420 236964 16268
rect 237020 4676 237076 20104
rect 238588 17668 238644 20104
rect 238588 17602 238644 17612
rect 238700 20076 240128 20132
rect 240380 20076 241696 20132
rect 241948 20076 243264 20132
rect 243628 20076 244832 20132
rect 237020 4610 237076 4620
rect 238588 16212 238644 16222
rect 237804 480 237972 532
rect 237804 476 238168 480
rect 237804 420 237860 476
rect 236908 364 237860 420
rect 237916 392 238168 476
rect 237944 -960 238168 392
rect 238588 420 238644 16156
rect 238700 4452 238756 20076
rect 238700 4386 238756 4396
rect 240268 16436 240324 16446
rect 239708 480 239876 532
rect 239708 476 240072 480
rect 239708 420 239764 476
rect 238588 364 239764 420
rect 239820 392 240072 476
rect 239848 -960 240072 392
rect 240268 420 240324 16380
rect 240380 4564 240436 20076
rect 241948 6132 242004 20076
rect 241948 6066 242004 6076
rect 240380 4498 240436 4508
rect 243628 4116 243684 20076
rect 246428 16100 246484 20104
rect 246428 16034 246484 16044
rect 247100 20076 247968 20132
rect 248668 20076 249536 20132
rect 250348 20076 251104 20132
rect 246988 14644 247044 14654
rect 245532 14532 245588 14542
rect 243628 4050 243684 4060
rect 243740 14308 243796 14318
rect 241612 480 241780 532
rect 243740 480 243796 14252
rect 245532 480 245588 14476
rect 241612 476 241976 480
rect 241612 420 241668 476
rect 240268 364 241668 420
rect 241724 392 241976 476
rect 241752 -960 241976 392
rect 243656 -960 243880 480
rect 245532 392 245784 480
rect 245560 -960 245784 392
rect 246988 420 247044 14588
rect 247100 7588 247156 20076
rect 247100 7522 247156 7532
rect 248668 4340 248724 20076
rect 248668 4274 248724 4284
rect 248780 14420 248836 14430
rect 247324 480 247492 532
rect 247324 476 247688 480
rect 247324 420 247380 476
rect 246988 364 247380 420
rect 247436 392 247688 476
rect 247464 -960 247688 392
rect 248780 420 248836 14364
rect 250348 4788 250404 20076
rect 252028 14868 252084 14878
rect 250348 4722 250404 4732
rect 250460 14756 250516 14766
rect 249228 480 249396 532
rect 249228 476 249592 480
rect 249228 420 249284 476
rect 248780 364 249284 420
rect 249340 392 249592 476
rect 249368 -960 249592 392
rect 250460 420 250516 14700
rect 251132 480 251300 532
rect 251132 476 251496 480
rect 251132 420 251188 476
rect 250460 364 251188 420
rect 251244 392 251496 476
rect 251272 -960 251496 392
rect 252028 420 252084 14812
rect 252700 9268 252756 20104
rect 253820 20076 254240 20132
rect 255388 20076 255808 20132
rect 252700 9202 252756 9212
rect 253708 14980 253764 14990
rect 253036 480 253204 532
rect 253036 476 253400 480
rect 253036 420 253092 476
rect 252028 364 253092 420
rect 253148 392 253400 476
rect 253176 -960 253400 392
rect 253708 420 253764 14924
rect 253820 6020 253876 20076
rect 253820 5954 253876 5964
rect 255388 3892 255444 20076
rect 257404 16884 257460 20104
rect 258748 20076 258944 20132
rect 257404 16818 257460 16828
rect 257852 17668 257908 17678
rect 255388 3826 255444 3836
rect 257068 4676 257124 4686
rect 254940 480 255108 532
rect 257068 480 257124 4620
rect 257852 4228 257908 17612
rect 257852 4162 257908 4172
rect 258748 4004 258804 20076
rect 260540 17668 260596 20104
rect 260540 17602 260596 17612
rect 261212 16884 261268 16894
rect 261212 7812 261268 16828
rect 262108 15988 262164 20104
rect 262108 15922 262164 15932
rect 262668 20076 263648 20132
rect 263788 20076 265216 20132
rect 265468 20076 266784 20132
rect 267260 20076 268352 20132
rect 268828 20076 269920 20132
rect 262668 8428 262724 20076
rect 261212 7746 261268 7756
rect 262108 8372 262724 8428
rect 262108 5908 262164 8372
rect 262108 5842 262164 5852
rect 262668 4564 262724 4574
rect 260764 4452 260820 4462
rect 258748 3938 258804 3948
rect 258860 4228 258916 4238
rect 258860 480 258916 4172
rect 260764 480 260820 4396
rect 262668 480 262724 4508
rect 263788 4564 263844 20076
rect 265468 7700 265524 20076
rect 265468 7634 265524 7644
rect 267148 16100 267204 16110
rect 263788 4498 263844 4508
rect 264572 6132 264628 6142
rect 264572 480 264628 6076
rect 266476 4116 266532 4126
rect 266476 480 266532 4060
rect 254940 476 255304 480
rect 254940 420 254996 476
rect 253708 364 254996 420
rect 255052 392 255304 476
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258860 392 259112 480
rect 260764 392 261016 480
rect 262668 392 262920 480
rect 264572 392 264824 480
rect 266476 392 266728 480
rect 258888 -960 259112 392
rect 260792 -960 261016 392
rect 262696 -960 262920 392
rect 264600 -960 264824 392
rect 266504 -960 266728 392
rect 267148 420 267204 16044
rect 267260 4676 267316 20076
rect 267260 4610 267316 4620
rect 268828 4228 268884 20076
rect 271516 16100 271572 20104
rect 273084 17220 273140 20104
rect 273084 17154 273140 17164
rect 273868 20076 274624 20132
rect 271516 16034 271572 16044
rect 268828 4162 268884 4172
rect 270284 7588 270340 7598
rect 268268 480 268436 532
rect 270284 480 270340 7532
rect 273868 4452 273924 20076
rect 276220 17892 276276 20104
rect 276220 17826 276276 17836
rect 275436 17220 275492 17230
rect 275436 14420 275492 17164
rect 275436 14354 275492 14364
rect 277788 12740 277844 20104
rect 277788 12674 277844 12684
rect 278908 20076 279328 20132
rect 280588 20076 280896 20132
rect 282268 20076 282464 20132
rect 283948 20076 284032 20132
rect 275996 9268 276052 9278
rect 273868 4386 273924 4396
rect 274092 4788 274148 4798
rect 272188 4340 272244 4350
rect 272188 480 272244 4284
rect 274092 480 274148 4732
rect 275996 480 276052 9212
rect 277900 6020 277956 6030
rect 277900 480 277956 5964
rect 278908 5012 278964 20076
rect 280588 7588 280644 20076
rect 280588 7522 280644 7532
rect 281708 7812 281764 7822
rect 278908 4946 278964 4956
rect 279804 4004 279860 4014
rect 279804 480 279860 3948
rect 281708 480 281764 7756
rect 282268 4900 282324 20076
rect 283948 6020 284004 20076
rect 285516 17668 285572 17678
rect 285516 16660 285572 17612
rect 285628 16884 285684 20104
rect 285628 16818 285684 16828
rect 285740 20076 287168 20132
rect 285516 16604 285684 16660
rect 283948 5954 284004 5964
rect 282268 4834 282324 4844
rect 283612 4116 283668 4126
rect 283612 480 283668 4060
rect 285628 480 285684 16604
rect 285740 4340 285796 20076
rect 288764 17668 288820 20104
rect 288764 17602 288820 17612
rect 289772 17892 289828 17902
rect 288764 16884 288820 16894
rect 285740 4274 285796 4284
rect 287420 15988 287476 15998
rect 287420 480 287476 15932
rect 288764 15988 288820 16828
rect 288764 15922 288820 15932
rect 289772 7924 289828 17836
rect 290332 17780 290388 20104
rect 291900 17892 291956 20104
rect 291900 17826 291956 17836
rect 292348 20076 293440 20132
rect 290332 17714 290388 17724
rect 289772 7858 289828 7868
rect 289324 5908 289380 5918
rect 289324 480 289380 5852
rect 292348 5908 292404 20076
rect 295036 16884 295092 20104
rect 295036 16818 295092 16828
rect 296492 16884 296548 16894
rect 296492 7812 296548 16828
rect 296604 14308 296660 20104
rect 297500 20076 298144 20132
rect 296604 14242 296660 14252
rect 297388 16100 297444 16110
rect 296492 7746 296548 7756
rect 292348 5842 292404 5852
rect 293132 7700 293188 7710
rect 291228 4564 291284 4574
rect 291228 480 291284 4508
rect 293132 480 293188 7644
rect 295036 4676 295092 4686
rect 295036 480 295092 4620
rect 296940 4228 296996 4238
rect 296940 480 296996 4172
rect 268268 476 268632 480
rect 268268 420 268324 476
rect 267148 364 268324 420
rect 268380 392 268632 476
rect 270284 392 270536 480
rect 272188 392 272440 480
rect 274092 392 274344 480
rect 275996 392 276248 480
rect 277900 392 278152 480
rect 279804 392 280056 480
rect 281708 392 281960 480
rect 283612 392 283864 480
rect 268408 -960 268632 392
rect 270312 -960 270536 392
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 276024 -960 276248 392
rect 277928 -960 278152 392
rect 279832 -960 280056 392
rect 281736 -960 281960 392
rect 283640 -960 283864 392
rect 285544 -960 285768 480
rect 287420 392 287672 480
rect 289324 392 289576 480
rect 291228 392 291480 480
rect 293132 392 293384 480
rect 295036 392 295288 480
rect 296940 392 297192 480
rect 287448 -960 287672 392
rect 289352 -960 289576 392
rect 291256 -960 291480 392
rect 293160 -960 293384 392
rect 295064 -960 295288 392
rect 296968 -960 297192 392
rect 297388 420 297444 16044
rect 297500 4788 297556 20076
rect 299740 10948 299796 20104
rect 299740 10882 299796 10892
rect 300748 14420 300804 14430
rect 297500 4722 297556 4732
rect 298732 480 298900 532
rect 300748 480 300804 14364
rect 301308 12628 301364 20104
rect 301308 12562 301364 12572
rect 302428 20076 302848 20132
rect 304108 20076 304416 20132
rect 302428 4228 302484 20076
rect 304108 7700 304164 20076
rect 305788 12740 305844 12750
rect 304108 7634 304164 7644
rect 304556 7924 304612 7934
rect 302428 4162 302484 4172
rect 302652 4452 302708 4462
rect 302652 480 302708 4396
rect 304556 480 304612 7868
rect 298732 476 299096 480
rect 298732 420 298788 476
rect 297388 364 298788 420
rect 298844 392 299096 476
rect 300748 392 301000 480
rect 302652 392 302904 480
rect 304556 392 304808 480
rect 298872 -960 299096 392
rect 300776 -960 301000 392
rect 302680 -960 302904 392
rect 304584 -960 304808 392
rect 305788 420 305844 12684
rect 306012 9268 306068 20104
rect 307468 20076 307552 20132
rect 306908 17892 306964 17902
rect 306908 12740 306964 17836
rect 306908 12674 306964 12684
rect 306012 9202 306068 9212
rect 307468 4676 307524 20076
rect 308252 17668 308308 17678
rect 307468 4610 307524 4620
rect 307580 7588 307636 7598
rect 307580 4564 307636 7532
rect 308252 6244 308308 17612
rect 309148 17668 309204 20104
rect 309148 17602 309204 17612
rect 310716 16884 310772 20104
rect 310716 16818 310772 16828
rect 310828 20076 312256 20132
rect 308252 6178 308308 6188
rect 307580 4498 307636 4508
rect 308364 5012 308420 5022
rect 306348 480 306516 532
rect 308364 480 308420 4956
rect 310268 4564 310324 4574
rect 310268 480 310324 4508
rect 310828 4564 310884 20076
rect 312396 16884 312452 16894
rect 312396 11060 312452 16828
rect 313852 16884 313908 20104
rect 313852 16818 313908 16828
rect 314972 17780 315028 17790
rect 312396 10994 312452 11004
rect 314972 6804 315028 17724
rect 315420 16212 315476 20104
rect 316988 17780 317044 20104
rect 316988 17714 317044 17724
rect 317548 20076 318528 20132
rect 315420 16146 315476 16156
rect 316652 16884 316708 16894
rect 314972 6738 315028 6748
rect 315980 15988 316036 15998
rect 314188 6020 314244 6030
rect 310828 4498 310884 4508
rect 312172 4900 312228 4910
rect 312172 480 312228 4844
rect 314188 480 314244 5964
rect 315980 480 316036 15932
rect 316652 14420 316708 16828
rect 316652 14354 316708 14364
rect 317548 6132 317604 20076
rect 320124 9380 320180 20104
rect 320124 9314 320180 9324
rect 320908 20076 321664 20132
rect 322700 20076 323232 20132
rect 324268 20076 324800 20132
rect 317548 6066 317604 6076
rect 319788 6244 319844 6254
rect 317884 4340 317940 4350
rect 317884 480 317940 4284
rect 319788 480 319844 6188
rect 320908 4452 320964 20076
rect 322588 12740 322644 12750
rect 320908 4386 320964 4396
rect 321692 6804 321748 6814
rect 321692 480 321748 6748
rect 306348 476 306712 480
rect 306348 420 306404 476
rect 305788 364 306404 420
rect 306460 392 306712 476
rect 308364 392 308616 480
rect 310268 392 310520 480
rect 312172 392 312424 480
rect 306488 -960 306712 392
rect 308392 -960 308616 392
rect 310296 -960 310520 392
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 315980 392 316232 480
rect 317884 392 318136 480
rect 319788 392 320040 480
rect 321692 392 321944 480
rect 316008 -960 316232 392
rect 317912 -960 318136 392
rect 319816 -960 320040 392
rect 321720 -960 321944 392
rect 322588 420 322644 12684
rect 322700 7588 322756 20076
rect 322700 7522 322756 7532
rect 324268 2548 324324 20076
rect 326396 17892 326452 20104
rect 326396 17826 326452 17836
rect 327628 20076 327936 20132
rect 327404 7812 327460 7822
rect 324268 2482 324324 2492
rect 325500 5908 325556 5918
rect 323484 480 323652 532
rect 325500 480 325556 5852
rect 327404 480 327460 7756
rect 327628 6020 327684 20076
rect 329532 15988 329588 20104
rect 329532 15922 329588 15932
rect 330988 20076 331072 20132
rect 327628 5954 327684 5964
rect 329308 14308 329364 14318
rect 329308 480 329364 14252
rect 330988 4340 331044 20076
rect 332668 16884 332724 20104
rect 332668 16818 332724 16828
rect 333116 10948 333172 10958
rect 330988 4274 331044 4284
rect 331212 4788 331268 4798
rect 331212 480 331268 4732
rect 333116 480 333172 10892
rect 334236 10948 334292 20104
rect 335804 18004 335860 20104
rect 335804 17938 335860 17948
rect 336812 17668 336868 17678
rect 335356 16884 335412 16894
rect 335356 14308 335412 16828
rect 335356 14242 335412 14252
rect 334236 10882 334292 10892
rect 334348 12628 334404 12638
rect 323484 476 323848 480
rect 323484 420 323540 476
rect 322588 364 323540 420
rect 323596 392 323848 476
rect 325500 392 325752 480
rect 327404 392 327656 480
rect 329308 392 329560 480
rect 331212 392 331464 480
rect 333116 392 333368 480
rect 323624 -960 323848 392
rect 325528 -960 325752 392
rect 327432 -960 327656 392
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 333144 -960 333368 392
rect 334348 420 334404 12572
rect 336812 6244 336868 17612
rect 337372 12740 337428 20104
rect 337372 12674 337428 12684
rect 337708 20076 338912 20132
rect 339388 20076 340480 20132
rect 341068 20076 342048 20132
rect 337708 7924 337764 20076
rect 337708 7858 337764 7868
rect 336812 6178 336868 6188
rect 338828 7700 338884 7710
rect 336924 4228 336980 4238
rect 334908 480 335076 532
rect 336924 480 336980 4172
rect 338828 480 338884 7644
rect 339388 4228 339444 20076
rect 339388 4162 339444 4172
rect 340732 9268 340788 9278
rect 340732 480 340788 9212
rect 341068 7812 341124 20076
rect 341068 7746 341124 7756
rect 343532 17780 343588 17790
rect 343532 5908 343588 17724
rect 343644 17332 343700 20104
rect 345240 20076 346052 20132
rect 343644 17266 343700 17276
rect 345996 16884 346052 20076
rect 346780 17780 346836 20104
rect 348376 20076 349300 20132
rect 346780 17714 346836 17724
rect 346892 17892 346948 17902
rect 345996 16828 346164 16884
rect 346108 12852 346164 16828
rect 346108 12786 346164 12796
rect 346444 11060 346500 11070
rect 343532 5842 343588 5852
rect 344540 6244 344596 6254
rect 342748 4676 342804 4686
rect 342748 480 342804 4620
rect 344540 480 344596 6188
rect 346444 480 346500 11004
rect 346892 6356 346948 17836
rect 349244 16884 349300 20076
rect 349244 16828 349524 16884
rect 349468 16100 349524 16828
rect 349468 16034 349524 16044
rect 346892 6290 346948 6300
rect 349468 14420 349524 14430
rect 348348 4564 348404 4574
rect 348348 480 348404 4508
rect 334908 476 335272 480
rect 334908 420 334964 476
rect 334348 364 334964 420
rect 335020 392 335272 476
rect 336924 392 337176 480
rect 338828 392 339080 480
rect 340732 392 340984 480
rect 335048 -960 335272 392
rect 336952 -960 337176 392
rect 338856 -960 339080 392
rect 340760 -960 340984 392
rect 342664 -960 342888 480
rect 344540 392 344792 480
rect 346444 392 346696 480
rect 348348 392 348600 480
rect 344568 -960 344792 392
rect 346472 -960 346696 392
rect 348376 -960 348600 392
rect 349468 420 349524 14364
rect 349916 11172 349972 20104
rect 351484 16884 351540 20104
rect 353052 17668 353108 20104
rect 354508 20076 354592 20132
rect 353052 17602 353108 17612
rect 353612 18004 353668 18014
rect 351484 16818 351540 16828
rect 352716 17332 352772 17342
rect 349916 11106 349972 11116
rect 351148 16212 351204 16222
rect 350140 480 350308 532
rect 350140 476 350504 480
rect 350140 420 350196 476
rect 349468 364 350196 420
rect 350252 392 350504 476
rect 350280 -960 350504 392
rect 351148 420 351204 16156
rect 352716 14420 352772 17276
rect 352716 14354 352772 14364
rect 353612 6244 353668 17948
rect 353612 6178 353668 6188
rect 354060 5908 354116 5918
rect 352044 480 352212 532
rect 354060 480 354116 5852
rect 354508 5908 354564 20076
rect 356188 18004 356244 20104
rect 356188 17938 356244 17948
rect 357756 9268 357812 20104
rect 359324 14644 359380 20104
rect 359324 14578 359380 14588
rect 360332 16884 360388 16894
rect 357756 9202 357812 9212
rect 357868 9380 357924 9390
rect 354508 5842 354564 5852
rect 355964 6132 356020 6142
rect 355964 480 356020 6076
rect 357868 480 357924 9324
rect 360332 8036 360388 16828
rect 360892 11060 360948 20104
rect 362460 12628 362516 20104
rect 364028 16884 364084 20104
rect 364028 16818 364084 16828
rect 365372 16884 365428 16894
rect 362460 12562 362516 12572
rect 360892 10994 360948 11004
rect 360332 7970 360388 7980
rect 361676 7588 361732 7598
rect 359772 4452 359828 4462
rect 359772 480 359828 4396
rect 361676 480 361732 7532
rect 365372 2996 365428 16828
rect 365596 9492 365652 20104
rect 367192 20076 367892 20132
rect 367836 18116 367892 20076
rect 367836 18060 368004 18116
rect 367948 15988 368004 18060
rect 368732 17892 368788 20104
rect 368732 17826 368788 17836
rect 369628 20076 370272 20132
rect 371420 20076 371840 20132
rect 367948 15922 368004 15932
rect 365596 9426 365652 9436
rect 367948 15764 368004 15774
rect 365372 2930 365428 2940
rect 365484 6356 365540 6366
rect 363580 2548 363636 2558
rect 363580 480 363636 2492
rect 365484 480 365540 6300
rect 367388 6020 367444 6030
rect 367388 480 367444 5964
rect 352044 476 352408 480
rect 352044 420 352100 476
rect 351148 364 352100 420
rect 352156 392 352408 476
rect 354060 392 354312 480
rect 355964 392 356216 480
rect 357868 392 358120 480
rect 359772 392 360024 480
rect 361676 392 361928 480
rect 363580 392 363832 480
rect 365484 392 365736 480
rect 367388 392 367640 480
rect 352184 -960 352408 392
rect 354088 -960 354312 392
rect 355992 -960 356216 392
rect 357896 -960 358120 392
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 363608 -960 363832 392
rect 365512 -960 365736 392
rect 367416 -960 367640 392
rect 367948 420 368004 15708
rect 369628 6020 369684 20076
rect 369628 5954 369684 5964
rect 371308 4340 371364 4350
rect 369180 480 369348 532
rect 371308 480 371364 4284
rect 371420 2660 371476 20076
rect 373436 16324 373492 20104
rect 375032 20076 375732 20132
rect 373436 16258 373492 16268
rect 374108 17780 374164 17790
rect 374108 14532 374164 17724
rect 374108 14466 374164 14476
rect 371420 2594 371476 2604
rect 373100 14308 373156 14318
rect 373100 480 373156 14252
rect 375676 10948 375732 20076
rect 376572 17780 376628 20104
rect 376572 17714 376628 17724
rect 377132 18004 377188 18014
rect 375676 10882 375732 10892
rect 375004 10836 375060 10846
rect 375004 480 375060 10780
rect 376908 6244 376964 6254
rect 376908 480 376964 6188
rect 377132 6132 377188 17948
rect 378140 14308 378196 20104
rect 379708 16884 379764 20104
rect 379708 16818 379764 16828
rect 380268 20076 381248 20132
rect 378140 14242 378196 14252
rect 377132 6066 377188 6076
rect 378028 12740 378084 12750
rect 369180 476 369544 480
rect 369180 420 369236 476
rect 367948 364 369236 420
rect 369292 392 369544 476
rect 369320 -960 369544 392
rect 371224 -960 371448 480
rect 373100 392 373352 480
rect 375004 392 375256 480
rect 376908 392 377160 480
rect 373128 -960 373352 392
rect 375032 -960 375256 392
rect 376936 -960 377160 392
rect 378028 420 378084 12684
rect 380268 8428 380324 20076
rect 382844 18004 382900 20104
rect 382844 17938 382900 17948
rect 383068 20076 384384 20132
rect 379708 8372 380324 8428
rect 379708 7700 379764 8372
rect 379708 7634 379764 7644
rect 380716 7924 380772 7934
rect 378700 480 378868 532
rect 380716 480 380772 7868
rect 383068 7588 383124 20076
rect 385980 18116 386036 20104
rect 385980 18050 386036 18060
rect 386428 20076 387520 20132
rect 388220 20076 389088 20132
rect 383516 16884 383572 16894
rect 383516 13076 383572 16828
rect 383516 13010 383572 13020
rect 383068 7522 383124 7532
rect 384524 7812 384580 7822
rect 382620 4228 382676 4238
rect 382620 480 382676 4172
rect 384524 480 384580 7756
rect 386428 2548 386484 20076
rect 387996 17668 388052 17678
rect 386428 2482 386484 2492
rect 386540 14420 386596 14430
rect 386540 480 386596 14364
rect 387996 14420 388052 17612
rect 387996 14354 388052 14364
rect 388108 12852 388164 12862
rect 388108 4228 388164 12796
rect 388220 7924 388276 20076
rect 388892 17780 388948 17790
rect 388892 12964 388948 17724
rect 388892 12898 388948 12908
rect 389788 14532 389844 14542
rect 388220 7858 388276 7868
rect 388108 4172 388388 4228
rect 388332 480 388388 4172
rect 378700 476 379064 480
rect 378700 420 378756 476
rect 378028 364 378756 420
rect 378812 392 379064 476
rect 380716 392 380968 480
rect 382620 392 382872 480
rect 384524 392 384776 480
rect 378840 -960 379064 392
rect 380744 -960 380968 392
rect 382648 -960 382872 392
rect 384552 -960 384776 392
rect 386456 -960 386680 480
rect 388332 392 388584 480
rect 388360 -960 388584 392
rect 389788 420 389844 14476
rect 390684 14532 390740 20104
rect 392252 16212 392308 20104
rect 392252 16146 392308 16156
rect 393148 20076 393792 20132
rect 390684 14466 390740 14476
rect 391468 16100 391524 16110
rect 390124 480 390292 532
rect 390124 476 390488 480
rect 390124 420 390180 476
rect 389788 364 390180 420
rect 390236 392 390488 476
rect 390264 -960 390488 392
rect 391468 420 391524 16044
rect 393148 6356 393204 20076
rect 393148 6290 393204 6300
rect 394044 11172 394100 11182
rect 392028 480 392196 532
rect 394044 480 394100 11116
rect 395388 9380 395444 20104
rect 395388 9314 395444 9324
rect 396508 14420 396564 14430
rect 395948 8036 396004 8046
rect 395948 480 396004 7980
rect 392028 476 392392 480
rect 392028 420 392084 476
rect 391468 364 392084 420
rect 392140 392 392392 476
rect 394044 392 394296 480
rect 395948 392 396200 480
rect 392168 -960 392392 392
rect 394072 -960 394296 392
rect 395976 -960 396200 392
rect 396508 420 396564 14364
rect 396956 12852 397012 20104
rect 398524 17780 398580 20104
rect 398524 17714 398580 17724
rect 400092 16100 400148 20104
rect 400092 16034 400148 16044
rect 400652 18004 400708 18014
rect 396956 12786 397012 12796
rect 400652 6468 400708 17948
rect 401660 17668 401716 20104
rect 403228 18004 403284 20104
rect 403228 17938 403284 17948
rect 401660 17602 401716 17612
rect 404796 14420 404852 20104
rect 404796 14354 404852 14364
rect 404908 14644 404964 14654
rect 400652 6402 400708 6412
rect 403564 9268 403620 9278
rect 401660 6132 401716 6142
rect 399868 5908 399924 5918
rect 397740 480 397908 532
rect 399868 480 399924 5852
rect 401660 480 401716 6076
rect 403564 480 403620 9212
rect 397740 476 398104 480
rect 397740 420 397796 476
rect 396508 364 397796 420
rect 397852 392 398104 476
rect 397880 -960 398104 392
rect 399784 -960 400008 480
rect 401660 392 401912 480
rect 403564 392 403816 480
rect 401688 -960 401912 392
rect 403592 -960 403816 392
rect 404908 420 404964 14588
rect 406364 9268 406420 20104
rect 407932 18228 407988 20104
rect 407932 18162 407988 18172
rect 407596 18116 407652 18126
rect 406364 9202 406420 9212
rect 407372 11060 407428 11070
rect 405356 480 405524 532
rect 407372 480 407428 11004
rect 407596 11060 407652 18060
rect 409500 12740 409556 20104
rect 409500 12674 409556 12684
rect 409948 20076 411040 20132
rect 407596 10994 407652 11004
rect 408268 12628 408324 12638
rect 405356 476 405720 480
rect 405356 420 405412 476
rect 404908 364 405412 420
rect 405468 392 405720 476
rect 407372 392 407624 480
rect 405496 -960 405720 392
rect 407400 -960 407624 392
rect 408268 420 408324 12572
rect 409948 2772 410004 20076
rect 412076 18228 412132 18238
rect 412076 9604 412132 18172
rect 412636 11396 412692 20104
rect 412636 11330 412692 11340
rect 413308 20076 414176 20132
rect 412076 9538 412132 9548
rect 413084 9492 413140 9502
rect 409948 2706 410004 2716
rect 411180 2996 411236 3006
rect 409164 480 409332 532
rect 411180 480 411236 2940
rect 413084 480 413140 9436
rect 413308 5908 413364 20076
rect 413308 5842 413364 5852
rect 414092 17892 414148 17902
rect 414092 5460 414148 17836
rect 415772 16884 415828 20104
rect 417368 20076 418292 20132
rect 418236 16884 418292 20076
rect 418236 16828 418404 16884
rect 415772 16818 415828 16828
rect 414092 5394 414148 5404
rect 414988 15988 415044 15998
rect 414988 480 415044 15932
rect 418348 15988 418404 16828
rect 418348 15922 418404 15932
rect 418908 11284 418964 20104
rect 418908 11218 418964 11228
rect 419132 16884 419188 16894
rect 419132 6244 419188 16828
rect 420476 16884 420532 20104
rect 420476 16818 420532 16828
rect 419132 6178 419188 6188
rect 421708 16324 421764 16334
rect 418796 6020 418852 6030
rect 416892 5460 416948 5470
rect 416892 480 416948 5404
rect 418796 480 418852 5964
rect 420700 2660 420756 2670
rect 420700 480 420756 2604
rect 409164 476 409528 480
rect 409164 420 409220 476
rect 408268 364 409220 420
rect 409276 392 409528 476
rect 411180 392 411432 480
rect 413084 392 413336 480
rect 414988 392 415240 480
rect 416892 392 417144 480
rect 418796 392 419048 480
rect 420700 392 420952 480
rect 409304 -960 409528 392
rect 411208 -960 411432 392
rect 413112 -960 413336 392
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418824 -960 419048 392
rect 420728 -960 420952 392
rect 421708 420 421764 16268
rect 422044 14756 422100 20104
rect 422044 14690 422100 14700
rect 423612 12628 423668 20104
rect 423612 12562 423668 12572
rect 425068 20076 425152 20132
rect 424508 10948 424564 10958
rect 422492 480 422660 532
rect 424508 480 424564 10892
rect 422492 476 422856 480
rect 422492 420 422548 476
rect 421708 364 422548 420
rect 422604 392 422856 476
rect 424508 392 424760 480
rect 422632 -960 422856 392
rect 424536 -960 424760 392
rect 425068 84 425124 20076
rect 426748 17892 426804 20104
rect 426748 17826 426804 17836
rect 427532 20076 428288 20132
rect 427308 16884 427364 16894
rect 425180 12964 425236 12974
rect 425180 420 425236 12908
rect 427308 12964 427364 16828
rect 427308 12898 427364 12908
rect 427532 8428 427588 20076
rect 426748 8372 427588 8428
rect 428428 14308 428484 14318
rect 426748 2660 426804 8372
rect 426748 2594 426804 2604
rect 426300 480 426468 532
rect 428428 480 428484 14252
rect 429884 14308 429940 20104
rect 429884 14242 429940 14252
rect 430108 20076 431424 20132
rect 430108 6132 430164 20076
rect 430108 6066 430164 6076
rect 430220 13076 430276 13086
rect 430220 480 430276 13020
rect 433020 10948 433076 20104
rect 433020 10882 433076 10892
rect 433468 20076 434560 20132
rect 433468 7812 433524 20076
rect 436156 16884 436212 20104
rect 436156 16818 436212 16828
rect 436828 20076 437696 20132
rect 433468 7746 433524 7756
rect 432124 7700 432180 7710
rect 432124 480 432180 7644
rect 435932 7588 435988 7598
rect 434028 6468 434084 6478
rect 434028 480 434084 6412
rect 435932 480 435988 7532
rect 436828 7588 436884 20076
rect 439292 18228 439348 20104
rect 439292 18162 439348 18172
rect 440860 16436 440916 20104
rect 441868 20076 442400 20132
rect 440860 16370 440916 16380
rect 440972 16884 441028 16894
rect 436828 7522 436884 7532
rect 437836 11060 437892 11070
rect 437836 480 437892 11004
rect 440972 7924 441028 16828
rect 440972 7858 441028 7868
rect 441644 8036 441700 8046
rect 439740 2548 439796 2558
rect 439740 480 439796 2492
rect 441644 480 441700 7980
rect 441868 2548 441924 20076
rect 443996 18116 444052 20104
rect 443996 18050 444052 18060
rect 445340 20076 445536 20132
rect 446908 20076 447104 20132
rect 444332 18004 444388 18014
rect 441868 2482 441924 2492
rect 443548 14532 443604 14542
rect 443548 480 443604 14476
rect 444332 8036 444388 17948
rect 444332 7970 444388 7980
rect 445228 16212 445284 16222
rect 445228 4228 445284 16156
rect 445340 7700 445396 20076
rect 445340 7634 445396 7644
rect 446908 6018 446964 20076
rect 448700 18004 448756 20104
rect 448700 17938 448756 17948
rect 449372 17780 449428 17790
rect 449260 9380 449316 9390
rect 446908 5966 446910 6018
rect 446962 5966 446964 6018
rect 446908 5954 446964 5966
rect 447356 6356 447412 6366
rect 445228 4172 445508 4228
rect 445452 480 445508 4172
rect 447356 480 447412 6300
rect 448812 5908 448868 5918
rect 448812 5814 448868 5852
rect 449260 480 449316 9324
rect 449372 5124 449428 17724
rect 450268 17780 450324 20104
rect 450268 17714 450324 17724
rect 450380 18228 450436 18238
rect 450380 13076 450436 18172
rect 451836 14532 451892 20104
rect 453404 18228 453460 20104
rect 453404 18162 453460 18172
rect 454972 16324 455028 20104
rect 454972 16258 455028 16268
rect 456092 17668 456148 17678
rect 451836 14466 451892 14476
rect 453628 16100 453684 16110
rect 450380 13010 450436 13020
rect 449372 5058 449428 5068
rect 450268 12852 450324 12862
rect 426300 476 426664 480
rect 426300 420 426356 476
rect 425180 364 426356 420
rect 426412 392 426664 476
rect 425404 84 425460 94
rect 425068 28 425404 84
rect 425404 18 425460 28
rect 426440 -960 426664 392
rect 428344 -960 428568 480
rect 430220 392 430472 480
rect 432124 392 432376 480
rect 434028 392 434280 480
rect 435932 392 436184 480
rect 437836 392 438088 480
rect 439740 392 439992 480
rect 441644 392 441896 480
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 447356 392 447608 480
rect 449260 392 449512 480
rect 430248 -960 430472 392
rect 432152 -960 432376 392
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 437864 -960 438088 392
rect 439768 -960 439992 392
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 447384 -960 447608 392
rect 449288 -960 449512 392
rect 450268 420 450324 12796
rect 453068 5124 453124 5134
rect 451052 480 451220 532
rect 453068 480 453124 5068
rect 451052 476 451416 480
rect 451052 420 451108 476
rect 450268 364 451108 420
rect 451164 392 451416 476
rect 453068 392 453320 480
rect 451192 -960 451416 392
rect 453096 -960 453320 392
rect 453628 420 453684 16044
rect 456092 6692 456148 17612
rect 456540 16212 456596 20104
rect 458108 17668 458164 20104
rect 458108 17602 458164 17612
rect 459228 18004 459284 18014
rect 456540 16146 456596 16156
rect 459228 9492 459284 17948
rect 459676 14644 459732 20104
rect 459676 14578 459732 14588
rect 459228 9426 459284 9436
rect 460348 14420 460404 14430
rect 458780 8036 458836 8046
rect 456092 6626 456148 6636
rect 456988 6692 457044 6702
rect 456204 6020 456260 6030
rect 456204 5926 456260 5964
rect 456316 5908 456372 5918
rect 456316 5814 456372 5852
rect 454860 480 455028 532
rect 456988 480 457044 6636
rect 458780 480 458836 7980
rect 454860 476 455224 480
rect 454860 420 454916 476
rect 453628 364 454916 420
rect 454972 392 455224 476
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 458808 -960 459032 392
rect 460348 420 460404 14364
rect 461244 11060 461300 20104
rect 461244 10994 461300 11004
rect 462028 20076 462784 20132
rect 462028 4788 462084 20076
rect 464380 18004 464436 20104
rect 464380 17938 464436 17948
rect 464604 18228 464660 18238
rect 464492 9604 464548 9614
rect 462028 4722 462084 4732
rect 462588 9268 462644 9278
rect 460572 480 460740 532
rect 462588 480 462644 9212
rect 464492 480 464548 9548
rect 464604 2884 464660 18172
rect 464604 2818 464660 2828
rect 465388 12740 465444 12750
rect 460572 476 460936 480
rect 460572 420 460628 476
rect 460348 364 460628 420
rect 460684 392 460936 476
rect 462588 392 462840 480
rect 464492 392 464744 480
rect 460712 -960 460936 392
rect 462616 -960 462840 392
rect 464520 -960 464744 392
rect 465388 420 465444 12684
rect 465948 11172 466004 20104
rect 465948 11106 466004 11116
rect 467068 20076 467488 20132
rect 467068 4900 467124 20076
rect 467852 18116 467908 18126
rect 467852 6356 467908 18060
rect 469084 12852 469140 20104
rect 470652 18564 470708 20104
rect 470652 18498 470708 18508
rect 469084 12786 469140 12796
rect 467852 6290 467908 6300
rect 470204 11396 470260 11406
rect 467068 4834 467124 4844
rect 468300 2772 468356 2782
rect 466284 480 466452 532
rect 468300 480 468356 2716
rect 470204 480 470260 11340
rect 472108 5908 472164 5918
rect 472108 480 472164 5852
rect 472220 4676 472276 20104
rect 473788 16884 473844 20104
rect 475356 18116 475412 20104
rect 475356 18050 475412 18060
rect 475580 20076 476896 20132
rect 473788 16818 473844 16828
rect 475468 15988 475524 15998
rect 472220 4610 472276 4620
rect 474012 6244 474068 6254
rect 474012 480 474068 6188
rect 466284 476 466648 480
rect 466284 420 466340 476
rect 465388 364 466340 420
rect 466396 392 466648 476
rect 468300 392 468552 480
rect 470204 392 470456 480
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 466424 -960 466648 392
rect 468328 -960 468552 392
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475468 420 475524 15932
rect 475580 4564 475636 20076
rect 477932 17892 477988 17902
rect 475580 4498 475636 4508
rect 477820 11284 477876 11294
rect 475804 480 475972 532
rect 477820 480 477876 11228
rect 477932 6244 477988 17836
rect 478492 14420 478548 20104
rect 478492 14354 478548 14364
rect 477932 6178 477988 6188
rect 478828 12964 478884 12974
rect 475804 476 476168 480
rect 475804 420 475860 476
rect 475468 364 475860 420
rect 475916 392 476168 476
rect 477820 392 478072 480
rect 475944 -960 476168 392
rect 477848 -960 478072 392
rect 478828 420 478884 12908
rect 480060 9268 480116 20104
rect 481628 17892 481684 20104
rect 481628 17826 481684 17836
rect 480844 16884 480900 16894
rect 480060 9202 480116 9212
rect 480508 14756 480564 14766
rect 479612 480 479780 532
rect 479612 476 479976 480
rect 479612 420 479668 476
rect 478828 364 479668 420
rect 479724 392 479976 476
rect 479752 -960 479976 392
rect 480508 420 480564 14700
rect 480844 9380 480900 16828
rect 483196 12740 483252 20104
rect 483196 12674 483252 12684
rect 484652 18116 484708 18126
rect 480844 9314 480900 9324
rect 482188 12628 482244 12638
rect 481516 480 481684 532
rect 481516 476 481880 480
rect 481516 420 481572 476
rect 480508 364 481572 420
rect 481628 392 481880 476
rect 481656 -960 481880 392
rect 482188 420 482244 12572
rect 484652 2772 484708 18060
rect 484764 12628 484820 20104
rect 484764 12562 484820 12572
rect 485548 20076 486304 20132
rect 487228 20076 487872 20132
rect 485548 4452 485604 20076
rect 487228 5908 487284 20076
rect 489468 16884 489524 20104
rect 489468 16818 489524 16828
rect 490588 20076 491008 20132
rect 487228 5842 487284 5852
rect 487340 6244 487396 6254
rect 485548 4386 485604 4396
rect 484652 2706 484708 2716
rect 483420 480 483588 532
rect 485660 480 485828 532
rect 483420 476 483784 480
rect 483420 420 483476 476
rect 482188 364 483476 420
rect 483532 392 483784 476
rect 483560 -960 483784 392
rect 485464 476 485828 480
rect 485464 392 485716 476
rect 485464 -960 485688 392
rect 485772 84 485828 476
rect 487340 480 487396 6188
rect 490588 4340 490644 20076
rect 492604 18340 492660 20104
rect 492604 18274 492660 18284
rect 492156 16884 492212 16894
rect 492156 16100 492212 16828
rect 492156 16034 492212 16044
rect 490588 4274 490644 4284
rect 490700 14308 490756 14318
rect 489244 2660 489300 2670
rect 489244 480 489300 2604
rect 487340 392 487592 480
rect 489244 392 489496 480
rect 485772 18 485828 28
rect 487368 -960 487592 392
rect 489272 -960 489496 392
rect 490700 420 490756 14252
rect 494172 10836 494228 20104
rect 495740 18116 495796 20104
rect 495740 18050 495796 18060
rect 496412 17892 496468 17902
rect 494172 10770 494228 10780
rect 494956 10948 495012 10958
rect 493052 6132 493108 6142
rect 491036 480 491204 532
rect 493052 480 493108 6076
rect 494956 480 495012 10892
rect 496412 7812 496468 17836
rect 497308 15988 497364 20104
rect 498876 18228 498932 20104
rect 498876 18162 498932 18172
rect 498988 20076 500416 20132
rect 497308 15922 497364 15932
rect 498092 17668 498148 17678
rect 496412 7746 496468 7756
rect 496860 7924 496916 7934
rect 496860 480 496916 7868
rect 498092 7924 498148 17612
rect 498092 7858 498148 7868
rect 498764 8036 498820 8046
rect 498764 480 498820 7980
rect 498988 4228 499044 20076
rect 502012 17892 502068 20104
rect 503608 20076 503972 20132
rect 502012 17826 502068 17836
rect 503132 18004 503188 18014
rect 501452 17780 501508 17790
rect 498988 4162 499044 4172
rect 500668 7588 500724 7598
rect 500668 480 500724 7532
rect 501452 6244 501508 17724
rect 501452 6178 501508 6188
rect 502572 13076 502628 13086
rect 502572 480 502628 13020
rect 503132 6132 503188 17948
rect 503916 16884 503972 20076
rect 505148 17668 505204 20104
rect 519372 20020 519428 522620
rect 521612 362964 521668 534604
rect 523292 532980 523348 532990
rect 521612 362898 521668 362908
rect 522508 519426 522564 519438
rect 522508 519374 522510 519426
rect 522562 519374 522564 519426
rect 522508 20132 522564 519374
rect 523292 430164 523348 532924
rect 523292 430098 523348 430108
rect 526652 112644 526708 544348
rect 556892 541044 556948 541054
rect 545132 536228 545188 536238
rect 540092 534436 540148 534446
rect 535052 531300 535108 531310
rect 533372 526148 533428 526158
rect 526652 112578 526708 112588
rect 530908 522788 530964 522798
rect 522508 20066 522564 20076
rect 519372 19954 519428 19964
rect 505148 17602 505204 17612
rect 506492 18340 506548 18350
rect 503916 16828 504084 16884
rect 504028 14308 504084 16828
rect 504028 14242 504084 14252
rect 504140 16436 504196 16446
rect 504140 8428 504196 16380
rect 503132 6066 503188 6076
rect 504028 8372 504196 8428
rect 491036 476 491400 480
rect 491036 420 491092 476
rect 490700 364 491092 420
rect 491148 392 491400 476
rect 493052 392 493304 480
rect 494956 392 495208 480
rect 496860 392 497112 480
rect 498764 392 499016 480
rect 500668 392 500920 480
rect 502572 392 502824 480
rect 491176 -960 491400 392
rect 493080 -960 493304 392
rect 494984 -960 495208 392
rect 496888 -960 497112 392
rect 498792 -960 499016 392
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 504028 420 504084 8372
rect 506492 7588 506548 18284
rect 513212 18228 513268 18238
rect 506492 7522 506548 7532
rect 510188 7700 510244 7710
rect 508284 6356 508340 6366
rect 506380 2548 506436 2558
rect 504364 480 504532 532
rect 506380 480 506436 2492
rect 508284 480 508340 6300
rect 510188 480 510244 7644
rect 512092 6020 512148 6030
rect 512092 480 512148 5964
rect 513212 6020 513268 18172
rect 520828 16324 520884 16334
rect 517468 14532 517524 14542
rect 513212 5954 513268 5964
rect 514108 9492 514164 9502
rect 514108 480 514164 9436
rect 515900 6244 515956 6254
rect 515900 480 515956 6188
rect 504364 476 504728 480
rect 504364 420 504420 476
rect 504028 364 504420 420
rect 504476 392 504728 476
rect 506380 392 506632 480
rect 508284 392 508536 480
rect 510188 392 510440 480
rect 512092 392 512344 480
rect 504504 -960 504728 392
rect 506408 -960 506632 392
rect 508312 -960 508536 392
rect 510216 -960 510440 392
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515900 392 516152 480
rect 515928 -960 516152 392
rect 517468 420 517524 14476
rect 519708 2884 519764 2894
rect 517692 480 517860 532
rect 519708 480 519764 2828
rect 517692 476 518056 480
rect 517692 420 517748 476
rect 517468 364 517748 420
rect 517804 392 518056 476
rect 519708 392 519960 480
rect 517832 -960 518056 392
rect 519736 -960 519960 392
rect 520828 420 520884 16268
rect 522508 16212 522564 16222
rect 521500 480 521668 532
rect 521500 476 521864 480
rect 521500 420 521556 476
rect 520828 364 521556 420
rect 521612 392 521864 476
rect 521640 -960 521864 392
rect 522508 420 522564 16156
rect 525868 14644 525924 14654
rect 525420 7924 525476 7934
rect 523404 480 523572 532
rect 525420 480 525476 7868
rect 523404 476 523768 480
rect 523404 420 523460 476
rect 522508 364 523460 420
rect 523516 392 523768 476
rect 525420 392 525672 480
rect 523544 -960 523768 392
rect 525448 -960 525672 392
rect 525868 420 525924 14588
rect 529228 11060 529284 11070
rect 527212 480 527380 532
rect 529228 480 529284 11004
rect 530908 8484 530964 522732
rect 533372 270564 533428 526092
rect 535052 468804 535108 531244
rect 538412 530964 538468 530974
rect 536732 529732 536788 529742
rect 536732 509124 536788 529676
rect 536732 509058 536788 509068
rect 535052 468738 535108 468748
rect 533372 270498 533428 270508
rect 538412 151284 538468 530908
rect 540092 191604 540148 534380
rect 541772 519428 541828 519438
rect 541772 231924 541828 519372
rect 545132 349524 545188 536172
rect 553532 536004 553588 536014
rect 548492 532868 548548 532878
rect 548492 389844 548548 532812
rect 550172 524580 550228 524590
rect 550172 416724 550228 524524
rect 551852 521220 551908 521230
rect 551852 495684 551908 521164
rect 551852 495618 551908 495628
rect 550172 416658 550228 416668
rect 548492 389778 548548 389788
rect 545132 349458 545188 349468
rect 541772 231858 541828 231868
rect 540092 191538 540148 191548
rect 538412 151218 538468 151228
rect 553532 58884 553588 535948
rect 555212 525924 555268 525934
rect 555212 99204 555268 525868
rect 556892 310884 556948 540988
rect 560252 539588 560308 539598
rect 556892 310818 556948 310828
rect 558572 539476 558628 539486
rect 558572 257124 558628 539420
rect 560252 297444 560308 539532
rect 563612 536116 563668 536126
rect 563612 336084 563668 536060
rect 566972 529508 567028 529518
rect 566972 455364 567028 529452
rect 566972 455298 567028 455308
rect 563612 336018 563668 336028
rect 560252 297378 560308 297388
rect 558572 257058 558628 257068
rect 568652 137844 568708 552860
rect 570332 551236 570388 551246
rect 570332 178164 570388 551180
rect 580412 539364 580468 539374
rect 575372 537908 575428 537918
rect 575372 376404 575428 537852
rect 575372 376338 575428 376348
rect 580412 218596 580468 539308
rect 590492 528052 590548 528062
rect 589596 524468 589652 524478
rect 589596 522788 589652 524412
rect 589596 522722 589652 522732
rect 590492 324548 590548 527996
rect 590604 523460 590660 588588
rect 593068 552804 593124 552814
rect 590604 523394 590660 523404
rect 590828 548996 590884 549006
rect 590828 523348 590884 548940
rect 590828 523282 590884 523292
rect 590492 324482 590548 324492
rect 580412 218530 580468 218540
rect 570332 178098 570388 178108
rect 568652 137778 568708 137788
rect 555212 99138 555268 99148
rect 553532 58818 553588 58828
rect 593068 33796 593124 552748
rect 593516 551124 593572 551134
rect 593404 546084 593460 546094
rect 593180 542836 593236 542846
rect 593180 483140 593236 542780
rect 593180 483074 593236 483084
rect 593292 529284 593348 529294
rect 593068 33730 593124 33740
rect 593292 20580 593348 529228
rect 593404 47012 593460 546028
rect 593516 73444 593572 551068
rect 593852 549444 593908 549454
rect 593628 524244 593684 524254
rect 593628 86660 593684 524188
rect 593740 520884 593796 520894
rect 593740 126308 593796 520828
rect 593852 165956 593908 549388
rect 594412 541268 594468 541278
rect 594188 527604 594244 527614
rect 593964 520996 594020 521006
rect 593964 205604 594020 520940
rect 594076 519316 594132 519326
rect 594076 245252 594132 519260
rect 594188 284900 594244 527548
rect 594300 526036 594356 526046
rect 594300 403844 594356 525980
rect 594412 443492 594468 541212
rect 594412 443426 594468 443436
rect 594524 519204 594580 519214
rect 594300 403778 594356 403788
rect 594188 284834 594244 284844
rect 594076 245186 594132 245196
rect 593964 205538 594020 205548
rect 593852 165890 593908 165900
rect 593740 126242 593796 126252
rect 593628 86594 593684 86604
rect 593516 73378 593572 73388
rect 593404 46946 593460 46956
rect 593292 20514 593348 20524
rect 539308 18564 539364 18574
rect 531468 18116 531524 18126
rect 531468 11060 531524 18060
rect 537628 12852 537684 12862
rect 531468 10994 531524 11004
rect 534940 11172 534996 11182
rect 530908 8418 530964 8428
rect 533036 6132 533092 6142
rect 531132 4788 531188 4798
rect 531132 480 531188 4732
rect 533036 480 533092 6076
rect 534940 480 534996 11116
rect 536844 4900 536900 4910
rect 536844 480 536900 4844
rect 527212 476 527576 480
rect 527212 420 527268 476
rect 525868 364 527268 420
rect 527324 392 527576 476
rect 529228 392 529480 480
rect 531132 392 531384 480
rect 533036 392 533288 480
rect 534940 392 535192 480
rect 536844 392 537096 480
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 -960 531384 392
rect 533064 -960 533288 392
rect 534968 -960 535192 392
rect 536872 -960 537096 392
rect 537628 420 537684 12796
rect 538636 480 538804 532
rect 538636 476 539000 480
rect 538636 420 538692 476
rect 537628 364 538692 420
rect 538748 392 539000 476
rect 538776 -960 539000 392
rect 539308 420 539364 18508
rect 548492 17892 548548 17902
rect 544460 9380 544516 9390
rect 542668 4676 542724 4686
rect 540540 480 540708 532
rect 542668 480 542724 4620
rect 544460 480 544516 9324
rect 548492 7700 548548 17836
rect 577052 17668 577108 17678
rect 562828 16100 562884 16110
rect 548492 7634 548548 7644
rect 549388 14420 549444 14430
rect 548268 4564 548324 4574
rect 546364 2772 546420 2782
rect 546364 480 546420 2716
rect 548268 480 548324 4508
rect 540540 476 540904 480
rect 540540 420 540596 476
rect 539308 364 540596 420
rect 540652 392 540904 476
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544460 392 544712 480
rect 546364 392 546616 480
rect 548268 392 548520 480
rect 544488 -960 544712 392
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 549388 420 549444 14364
rect 554428 12740 554484 12750
rect 552076 9268 552132 9278
rect 550060 480 550228 532
rect 552076 480 552132 9212
rect 553980 7812 554036 7822
rect 553980 480 554036 7756
rect 550060 476 550424 480
rect 550060 420 550116 476
rect 549388 364 550116 420
rect 550172 392 550424 476
rect 552076 392 552328 480
rect 553980 392 554232 480
rect 550200 -960 550424 392
rect 552104 -960 552328 392
rect 554008 -960 554232 392
rect 554428 420 554484 12684
rect 557788 12628 557844 12638
rect 555772 480 555940 532
rect 557788 480 557844 12572
rect 561036 5908 561092 5918
rect 561036 5012 561092 5852
rect 561036 4956 561204 5012
rect 559692 4452 559748 4462
rect 559692 480 559748 4396
rect 555772 476 556136 480
rect 555772 420 555828 476
rect 554428 364 555828 420
rect 555884 392 556136 476
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561148 420 561204 4956
rect 561484 480 561652 532
rect 561484 476 561848 480
rect 561484 420 561540 476
rect 561148 364 561540 420
rect 561596 392 561848 476
rect 561624 -960 561848 392
rect 562828 420 562884 16044
rect 573020 15988 573076 15998
rect 571228 11060 571284 11070
rect 569212 10948 569268 10958
rect 567308 7588 567364 7598
rect 565404 4340 565460 4350
rect 563388 480 563556 532
rect 565404 480 565460 4284
rect 567308 480 567364 7532
rect 569212 480 569268 10892
rect 571228 480 571284 11004
rect 573020 480 573076 15932
rect 574924 6020 574980 6030
rect 574924 480 574980 5964
rect 577052 4788 577108 17612
rect 581308 14308 581364 14318
rect 577052 4722 577108 4732
rect 580636 7700 580692 7710
rect 576828 4228 576884 4238
rect 576828 480 576884 4172
rect 580636 480 580692 7644
rect 563388 476 563752 480
rect 563388 420 563444 476
rect 562828 364 563444 420
rect 563500 392 563752 476
rect 565404 392 565656 480
rect 567308 392 567560 480
rect 569212 392 569464 480
rect 563528 -960 563752 392
rect 565432 -960 565656 392
rect 567336 -960 567560 392
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 574924 392 575176 480
rect 576828 392 577080 480
rect 573048 -960 573272 392
rect 574952 -960 575176 392
rect 576856 -960 577080 392
rect 578760 -960 578984 480
rect 580636 392 580888 480
rect 580664 -960 580888 392
rect 581308 420 581364 14252
rect 594524 7364 594580 519148
rect 594524 7298 594580 7308
rect 584444 4788 584500 4798
rect 582428 480 582596 532
rect 584444 480 584500 4732
rect 582428 476 582792 480
rect 582428 420 582484 476
rect 581308 364 582484 420
rect 582540 392 582792 476
rect 584444 392 584696 480
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 31948 577052 32004 577108
rect 53788 560252 53844 560308
rect 10108 556892 10164 556948
rect 5852 556108 5908 556164
rect 2492 547708 2548 547764
rect 140 532588 196 532644
rect 28 521052 84 521108
rect 140 220556 196 220612
rect 28 79436 84 79492
rect 2716 534492 2772 534548
rect 2604 527660 2660 527716
rect 5068 524636 5124 524692
rect 5068 516796 5124 516852
rect 2716 403900 2772 403956
rect 2604 305116 2660 305172
rect 17724 554428 17780 554484
rect 12572 547820 12628 547876
rect 9436 542892 9492 542948
rect 9212 542668 9268 542724
rect 5964 537628 6020 537684
rect 6076 519484 6132 519540
rect 6076 262780 6132 262836
rect 5964 192220 6020 192276
rect 5852 107436 5908 107492
rect 9324 529564 9380 529620
rect 9324 418012 9380 418068
rect 10892 541100 10948 541156
rect 9548 521276 9604 521332
rect 9548 502684 9604 502740
rect 9436 333340 9492 333396
rect 11004 537740 11060 537796
rect 11116 531132 11172 531188
rect 11116 389676 11172 389732
rect 11004 276892 11060 276948
rect 10892 248556 10948 248612
rect 15932 546140 15988 546196
rect 14476 539644 14532 539700
rect 14364 532700 14420 532756
rect 12796 527884 12852 527940
rect 12684 526204 12740 526260
rect 12796 445228 12852 445284
rect 14252 522508 14308 522564
rect 12684 346108 12740 346164
rect 12572 120988 12628 121044
rect 9212 93436 9268 93492
rect 14700 536284 14756 536340
rect 14588 522620 14644 522676
rect 14700 487228 14756 487284
rect 14588 473788 14644 473844
rect 14476 361340 14532 361396
rect 14364 176428 14420 176484
rect 17612 531020 17668 531076
rect 16156 526316 16212 526372
rect 16044 524300 16100 524356
rect 16156 431900 16212 431956
rect 16044 290780 16100 290836
rect 70588 552860 70644 552916
rect 26908 552748 26964 552804
rect 19292 549500 19348 549556
rect 17836 537964 17892 538020
rect 17836 317548 17892 317604
rect 17724 233548 17780 233604
rect 17612 204988 17668 205044
rect 19404 544572 19460 544628
rect 19516 527772 19572 527828
rect 40348 551068 40404 551124
rect 35308 546028 35364 546084
rect 32060 529228 32116 529284
rect 53788 544348 53844 544404
rect 44268 535948 44324 536004
rect 50092 524188 50148 524244
rect 66108 530908 66164 530964
rect 58492 525868 58548 525924
rect 63196 520828 63252 520884
rect 99148 570332 99204 570388
rect 77308 550172 77364 550228
rect 84028 551180 84084 551236
rect 75628 549388 75684 549444
rect 79212 534380 79268 534436
rect 119308 540988 119364 541044
rect 109228 539420 109284 539476
rect 97468 539308 97524 539364
rect 88956 520940 89012 520996
rect 106876 526092 106932 526148
rect 115612 527548 115668 527604
rect 165676 590156 165732 590212
rect 167132 590156 167188 590212
rect 187740 590156 187796 590212
rect 188972 590156 189028 590212
rect 167132 568652 167188 568708
rect 188972 566972 189028 567028
rect 142828 546812 142884 546868
rect 206668 548492 206724 548548
rect 179788 542780 179844 542836
rect 166348 541212 166404 541268
rect 122668 539532 122724 539588
rect 149548 537852 149604 537908
rect 120988 523628 121044 523684
rect 131628 536172 131684 536228
rect 128716 523516 128772 523572
rect 136108 536060 136164 536116
rect 141260 534604 141316 534660
rect 144732 532812 144788 532868
rect 157948 532924 158004 532980
rect 154476 525980 154532 526036
rect 163660 524524 163716 524580
rect 171388 531244 171444 531300
rect 175308 529452 175364 529508
rect 208348 543452 208404 543508
rect 220892 593068 220948 593124
rect 215068 541772 215124 541828
rect 201628 534268 201684 534324
rect 184940 529676 184996 529732
rect 194236 524412 194292 524468
rect 189756 521164 189812 521220
rect 198156 523292 198212 523348
rect 211596 523404 211652 523460
rect 219884 523180 219940 523236
rect 220892 523180 220948 523236
rect 223468 555212 223524 555268
rect 228508 551852 228564 551908
rect 242732 593292 242788 593348
rect 234332 593180 234388 593236
rect 232652 574588 232708 574644
rect 232652 541772 232708 541828
rect 230188 523740 230244 523796
rect 231868 527996 231924 528052
rect 231868 523516 231924 523572
rect 233436 522732 233492 522788
rect 234332 522732 234388 522788
rect 237916 523516 237972 523572
rect 241836 522732 241892 522788
rect 253932 588812 253988 588868
rect 261212 590492 261268 590548
rect 253708 563612 253764 563668
rect 242732 522732 242788 522788
rect 245308 553532 245364 553588
rect 250348 541772 250404 541828
rect 259756 522732 259812 522788
rect 274652 578732 274708 578788
rect 267148 565292 267204 565348
rect 262108 561932 262164 561988
rect 261212 522732 261268 522788
rect 272748 522732 272804 522788
rect 283948 588812 284004 588868
rect 280588 572012 280644 572068
rect 274652 522732 274708 522788
rect 319228 578732 319284 578788
rect 335132 590604 335188 590660
rect 297388 572012 297444 572068
rect 332668 577052 332724 577108
rect 319228 570332 319284 570388
rect 305788 568652 305844 568708
rect 297388 566972 297444 567028
rect 288988 543452 289044 543508
rect 302428 546812 302484 546868
rect 294140 523740 294196 523796
rect 315868 550172 315924 550228
rect 324268 560252 324324 560308
rect 310828 523628 310884 523684
rect 327628 556892 327684 556948
rect 335132 565292 335188 565348
rect 337708 586348 337764 586404
rect 364028 590604 364084 590660
rect 365372 590604 365428 590660
rect 341068 561932 341124 561988
rect 346108 572908 346164 572964
rect 343532 561148 343588 561204
rect 341068 557788 341124 557844
rect 343532 548492 343588 548548
rect 386092 590492 386148 590548
rect 365372 553532 365428 553588
rect 349468 544460 349524 544516
rect 452284 590604 452340 590660
rect 430108 563612 430164 563668
rect 450268 554428 450324 554484
rect 408268 541772 408324 541828
rect 414988 542892 415044 542948
rect 411628 539644 411684 539700
rect 371868 536284 371924 536340
rect 359660 529340 359716 529396
rect 354508 524636 354564 524692
rect 367948 522620 368004 522676
rect 363244 521276 363300 521332
rect 398188 534492 398244 534548
rect 393708 531132 393764 531188
rect 389788 529564 389844 529620
rect 385084 527884 385140 527940
rect 381500 526316 381556 526372
rect 403340 527772 403396 527828
rect 406924 526204 406980 526260
rect 441868 541100 441924 541156
rect 425068 537964 425124 538020
rect 436828 537740 436884 537796
rect 420028 527660 420084 527716
rect 428764 524300 428820 524356
rect 472108 546140 472164 546196
rect 468748 544572 468804 544628
rect 463708 537628 463764 537684
rect 447020 532588 447076 532644
rect 459228 532700 459284 532756
rect 455308 531020 455364 531076
rect 496412 593292 496468 593348
rect 518476 593180 518532 593236
rect 496412 590492 496468 590548
rect 490588 556108 490644 556164
rect 473788 523516 473844 523572
rect 477148 549500 477204 549556
rect 480508 547820 480564 547876
rect 485548 542668 485604 542724
rect 584668 593068 584724 593124
rect 562604 590492 562660 590548
rect 539308 555212 539364 555268
rect 590604 588588 590660 588644
rect 496412 551852 496468 551908
rect 568652 552860 568708 552916
rect 498988 547708 499044 547764
rect 494284 521052 494340 521108
rect 526652 544348 526708 544404
rect 521612 534604 521668 534660
rect 513100 522732 513156 522788
rect 508732 522620 508788 522676
rect 503020 522508 503076 522564
rect 519372 522620 519428 522676
rect 19628 519596 19684 519652
rect 377020 519596 377076 519652
rect 433804 519484 433860 519540
rect 93100 519372 93156 519428
rect 23212 519260 23268 519316
rect 101836 519260 101892 519316
rect 19628 458668 19684 458724
rect 19516 374668 19572 374724
rect 19404 162988 19460 163044
rect 19292 149660 19348 149716
rect 15932 134428 15988 134484
rect 14252 63868 14308 63924
rect 2492 51100 2548 51156
rect 4172 36764 4228 36820
rect 4956 22652 5012 22708
rect 4956 20076 5012 20132
rect 4172 19964 4228 20020
rect 32732 18284 32788 18340
rect 18508 17612 18564 17668
rect 15148 12572 15204 12628
rect 13356 10892 13412 10948
rect 11564 7532 11620 7588
rect 17276 4172 17332 4228
rect 30380 15932 30436 15988
rect 22988 5852 23044 5908
rect 21084 4284 21140 4340
rect 28700 4620 28756 4676
rect 24892 4508 24948 4564
rect 26796 4396 26852 4452
rect 31948 14252 32004 14308
rect 32732 5852 32788 5908
rect 33628 18060 33684 18116
rect 33740 7532 33796 7588
rect 35308 17948 35364 18004
rect 35644 10892 35700 10948
rect 36988 17836 37044 17892
rect 37212 12572 37268 12628
rect 38668 17724 38724 17780
rect 40348 17612 40404 17668
rect 40460 18172 40516 18228
rect 38780 4172 38836 4228
rect 43932 18284 43988 18340
rect 42028 4284 42084 4340
rect 43932 11004 43988 11060
rect 45388 4508 45444 4564
rect 45836 11564 45892 11620
rect 47068 4396 47124 4452
rect 47740 11228 47796 11284
rect 50428 15932 50484 15988
rect 52892 18060 52948 18116
rect 54460 17948 54516 18004
rect 56364 17836 56420 17892
rect 59164 18172 59220 18228
rect 57596 17724 57652 17780
rect 51324 14252 51380 14308
rect 60508 17612 60564 17668
rect 48748 4620 48804 4676
rect 49644 11452 49700 11508
rect 55356 11340 55412 11396
rect 51548 11116 51604 11172
rect 53452 10892 53508 10948
rect 57260 4284 57316 4340
rect 59164 4172 59220 4228
rect 60732 11004 60788 11060
rect 62188 17836 62244 17892
rect 62300 11564 62356 11620
rect 63868 17948 63924 18004
rect 63980 11228 64036 11284
rect 65548 17724 65604 17780
rect 65660 11452 65716 11508
rect 67228 18060 67284 18116
rect 67452 11116 67508 11172
rect 68908 10892 68964 10948
rect 69020 18172 69076 18228
rect 70588 11340 70644 11396
rect 72268 4284 72324 4340
rect 72380 13244 72436 13300
rect 74172 13132 74228 13188
rect 77980 17948 78036 18004
rect 76412 17836 76468 17892
rect 82684 18172 82740 18228
rect 81116 18060 81172 18116
rect 79884 17724 79940 17780
rect 74844 17612 74900 17668
rect 84252 13244 84308 13300
rect 85708 17724 85764 17780
rect 80668 13020 80724 13076
rect 77308 12796 77364 12852
rect 74284 4172 74340 4228
rect 75628 12684 75684 12740
rect 78988 12572 79044 12628
rect 82348 12908 82404 12964
rect 85820 13132 85876 13188
rect 89068 17948 89124 18004
rect 87388 12684 87444 12740
rect 87500 17612 87556 17668
rect 89180 12796 89236 12852
rect 90748 18172 90804 18228
rect 92428 13020 92484 13076
rect 92540 18284 92596 18340
rect 90972 12572 91028 12628
rect 94108 16940 94164 16996
rect 95788 17724 95844 17780
rect 97468 17612 97524 17668
rect 97692 18396 97748 18452
rect 94220 12908 94276 12964
rect 95900 16828 95956 16884
rect 101500 18284 101556 18340
rect 99932 18172 99988 18228
rect 98364 17948 98420 18004
rect 102732 18060 102788 18116
rect 100828 17612 100884 17668
rect 103516 16940 103572 16996
rect 104188 17948 104244 18004
rect 106204 18396 106260 18452
rect 104636 16828 104692 16884
rect 105868 18172 105924 18228
rect 109340 18060 109396 18116
rect 112588 18172 112644 18228
rect 110908 17948 110964 18004
rect 107772 17612 107828 17668
rect 110908 17724 110964 17780
rect 107660 16940 107716 16996
rect 109228 16828 109284 16884
rect 114268 17612 114324 17668
rect 114492 16940 114548 16996
rect 117628 17724 117684 17780
rect 119308 17612 119364 17668
rect 115948 16828 116004 16884
rect 116060 16940 116116 16996
rect 120988 16940 121044 16996
rect 117628 15036 117684 15092
rect 121884 15036 121940 15092
rect 122780 15036 122836 15092
rect 120988 14924 121044 14980
rect 119308 14700 119364 14756
rect 126924 15036 126980 15092
rect 125020 14924 125076 14980
rect 123452 14700 123508 14756
rect 126028 14812 126084 14868
rect 124348 14364 124404 14420
rect 129724 14812 129780 14868
rect 128156 14364 128212 14420
rect 131292 13356 131348 13412
rect 129388 13244 129444 13300
rect 132860 13356 132916 13412
rect 131404 13244 131460 13300
rect 132748 13244 132804 13300
rect 134428 13244 134484 13300
rect 134540 13356 134596 13412
rect 136108 13356 136164 13412
rect 137900 13244 137956 13300
rect 136108 12012 136164 12068
rect 138012 12012 138068 12068
rect 139468 13356 139524 13412
rect 141148 13356 141204 13412
rect 139580 13244 139636 13300
rect 144732 4620 144788 4676
rect 147868 4956 147924 5012
rect 146188 4284 146244 4340
rect 146524 4620 146580 4676
rect 148428 4284 148484 4340
rect 149548 4284 149604 4340
rect 150332 4956 150388 5012
rect 151228 4172 151284 4228
rect 152236 4284 152292 4340
rect 154588 4620 154644 4676
rect 152908 4284 152964 4340
rect 156044 4284 156100 4340
rect 154140 4172 154196 4228
rect 159628 4844 159684 4900
rect 158060 4732 158116 4788
rect 156268 4172 156324 4228
rect 157948 4620 158004 4676
rect 159852 4172 159908 4228
rect 161308 4172 161364 4228
rect 161756 4732 161812 4788
rect 162988 4284 163044 4340
rect 163660 4844 163716 4900
rect 168140 5964 168196 6020
rect 171388 6076 171444 6132
rect 169708 5852 169764 5908
rect 176428 6412 176484 6468
rect 174748 6188 174804 6244
rect 173068 5068 173124 5124
rect 175084 5964 175140 6020
rect 168028 4732 168084 4788
rect 173180 4732 173236 4788
rect 166348 4508 166404 4564
rect 171388 4508 171444 4564
rect 167468 4284 167524 4340
rect 164668 4060 164724 4116
rect 165564 4172 165620 4228
rect 169372 4060 169428 4116
rect 176988 5852 177044 5908
rect 178108 5740 178164 5796
rect 178892 6076 178948 6132
rect 181468 6076 181524 6132
rect 182700 6188 182756 6244
rect 179788 5852 179844 5908
rect 180796 5068 180852 5124
rect 183148 6188 183204 6244
rect 184604 6412 184660 6468
rect 186508 6300 186564 6356
rect 188188 5964 188244 6020
rect 188412 5852 188468 5908
rect 184828 5068 184884 5124
rect 186508 5740 186564 5796
rect 189868 4172 189924 4228
rect 190316 6076 190372 6132
rect 191660 6412 191716 6468
rect 191548 4284 191604 4340
rect 192220 6188 192276 6244
rect 194908 6188 194964 6244
rect 196028 6300 196084 6356
rect 193228 5964 193284 6020
rect 194124 5068 194180 5124
rect 196588 6300 196644 6356
rect 198268 6076 198324 6132
rect 197932 5852 197988 5908
rect 204092 11228 204148 11284
rect 207228 11564 207284 11620
rect 211932 11452 211988 11508
rect 210364 11340 210420 11396
rect 208796 11116 208852 11172
rect 205660 11004 205716 11060
rect 202524 10892 202580 10948
rect 199948 5852 200004 5908
rect 203644 6412 203700 6468
rect 201740 4284 201796 4340
rect 199948 4172 200004 4228
rect 209356 6300 209412 6356
rect 207452 6188 207508 6244
rect 205548 5964 205604 6020
rect 211260 6076 211316 6132
rect 213164 5852 213220 5908
rect 213388 5852 213444 5908
rect 215068 10892 215124 10948
rect 216636 16492 216692 16548
rect 218204 16044 218260 16100
rect 221340 16268 221396 16324
rect 224476 16380 224532 16436
rect 222908 16156 222964 16212
rect 219772 15932 219828 15988
rect 229180 14588 229236 14644
rect 227612 14476 227668 14532
rect 230748 14364 230804 14420
rect 231868 16492 231924 16548
rect 226044 14252 226100 14308
rect 220780 11564 220836 11620
rect 215180 5964 215236 6020
rect 216972 11228 217028 11284
rect 218876 11004 218932 11060
rect 226492 11452 226548 11508
rect 224588 11340 224644 11396
rect 222684 11116 222740 11172
rect 230300 5964 230356 6020
rect 228508 5852 228564 5908
rect 232316 14700 232372 14756
rect 233548 16044 233604 16100
rect 233884 14812 233940 14868
rect 235228 15932 235284 15988
rect 235452 14924 235508 14980
rect 236908 16268 236964 16324
rect 238588 17612 238644 17668
rect 237020 4620 237076 4676
rect 238588 16156 238644 16212
rect 238700 4396 238756 4452
rect 240268 16380 240324 16436
rect 241948 6076 242004 6132
rect 240380 4508 240436 4564
rect 246428 16044 246484 16100
rect 246988 14588 247044 14644
rect 245532 14476 245588 14532
rect 243628 4060 243684 4116
rect 243740 14252 243796 14308
rect 247100 7532 247156 7588
rect 248668 4284 248724 4340
rect 248780 14364 248836 14420
rect 252028 14812 252084 14868
rect 250348 4732 250404 4788
rect 250460 14700 250516 14756
rect 252700 9212 252756 9268
rect 253708 14924 253764 14980
rect 253820 5964 253876 6020
rect 257404 16828 257460 16884
rect 257852 17612 257908 17668
rect 255388 3836 255444 3892
rect 257068 4620 257124 4676
rect 257852 4172 257908 4228
rect 260540 17612 260596 17668
rect 261212 16828 261268 16884
rect 262108 15932 262164 15988
rect 261212 7756 261268 7812
rect 262108 5852 262164 5908
rect 262668 4508 262724 4564
rect 260764 4396 260820 4452
rect 258748 3948 258804 4004
rect 258860 4172 258916 4228
rect 265468 7644 265524 7700
rect 267148 16044 267204 16100
rect 263788 4508 263844 4564
rect 264572 6076 264628 6132
rect 266476 4060 266532 4116
rect 267260 4620 267316 4676
rect 273084 17164 273140 17220
rect 271516 16044 271572 16100
rect 268828 4172 268884 4228
rect 270284 7532 270340 7588
rect 276220 17836 276276 17892
rect 275436 17164 275492 17220
rect 275436 14364 275492 14420
rect 277788 12684 277844 12740
rect 275996 9212 276052 9268
rect 273868 4396 273924 4452
rect 274092 4732 274148 4788
rect 272188 4284 272244 4340
rect 277900 5964 277956 6020
rect 280588 7532 280644 7588
rect 281708 7756 281764 7812
rect 278908 4956 278964 5012
rect 279804 3948 279860 4004
rect 285516 17612 285572 17668
rect 285628 16828 285684 16884
rect 283948 5964 284004 6020
rect 282268 4844 282324 4900
rect 283612 4060 283668 4116
rect 288764 17612 288820 17668
rect 289772 17836 289828 17892
rect 288764 16828 288820 16884
rect 285740 4284 285796 4340
rect 287420 15932 287476 15988
rect 288764 15932 288820 15988
rect 291900 17836 291956 17892
rect 290332 17724 290388 17780
rect 289772 7868 289828 7924
rect 289324 5852 289380 5908
rect 295036 16828 295092 16884
rect 296492 16828 296548 16884
rect 296604 14252 296660 14308
rect 297388 16044 297444 16100
rect 296492 7756 296548 7812
rect 292348 5852 292404 5908
rect 293132 7644 293188 7700
rect 291228 4508 291284 4564
rect 295036 4620 295092 4676
rect 296940 4172 296996 4228
rect 299740 10892 299796 10948
rect 300748 14364 300804 14420
rect 297500 4732 297556 4788
rect 301308 12572 301364 12628
rect 305788 12684 305844 12740
rect 304108 7644 304164 7700
rect 304556 7868 304612 7924
rect 302428 4172 302484 4228
rect 302652 4396 302708 4452
rect 306908 17836 306964 17892
rect 306908 12684 306964 12740
rect 306012 9212 306068 9268
rect 308252 17612 308308 17668
rect 307468 4620 307524 4676
rect 307580 7532 307636 7588
rect 309148 17612 309204 17668
rect 310716 16828 310772 16884
rect 308252 6188 308308 6244
rect 307580 4508 307636 4564
rect 308364 4956 308420 5012
rect 310268 4508 310324 4564
rect 312396 16828 312452 16884
rect 313852 16828 313908 16884
rect 314972 17724 315028 17780
rect 312396 11004 312452 11060
rect 316988 17724 317044 17780
rect 315420 16156 315476 16212
rect 316652 16828 316708 16884
rect 314972 6748 315028 6804
rect 315980 15932 316036 15988
rect 314188 5964 314244 6020
rect 310828 4508 310884 4564
rect 312172 4844 312228 4900
rect 316652 14364 316708 14420
rect 320124 9324 320180 9380
rect 317548 6076 317604 6132
rect 319788 6188 319844 6244
rect 317884 4284 317940 4340
rect 322588 12684 322644 12740
rect 320908 4396 320964 4452
rect 321692 6748 321748 6804
rect 322700 7532 322756 7588
rect 326396 17836 326452 17892
rect 327404 7756 327460 7812
rect 324268 2492 324324 2548
rect 325500 5852 325556 5908
rect 329532 15932 329588 15988
rect 327628 5964 327684 6020
rect 329308 14252 329364 14308
rect 332668 16828 332724 16884
rect 333116 10892 333172 10948
rect 330988 4284 331044 4340
rect 331212 4732 331268 4788
rect 335804 17948 335860 18004
rect 336812 17612 336868 17668
rect 335356 16828 335412 16884
rect 335356 14252 335412 14308
rect 334236 10892 334292 10948
rect 334348 12572 334404 12628
rect 337372 12684 337428 12740
rect 337708 7868 337764 7924
rect 336812 6188 336868 6244
rect 338828 7644 338884 7700
rect 336924 4172 336980 4228
rect 339388 4172 339444 4228
rect 340732 9212 340788 9268
rect 341068 7756 341124 7812
rect 343532 17724 343588 17780
rect 343644 17276 343700 17332
rect 346780 17724 346836 17780
rect 346892 17836 346948 17892
rect 346108 12796 346164 12852
rect 346444 11004 346500 11060
rect 343532 5852 343588 5908
rect 344540 6188 344596 6244
rect 342748 4620 342804 4676
rect 349468 16044 349524 16100
rect 346892 6300 346948 6356
rect 349468 14364 349524 14420
rect 348348 4508 348404 4564
rect 353052 17612 353108 17668
rect 353612 17948 353668 18004
rect 351484 16828 351540 16884
rect 352716 17276 352772 17332
rect 349916 11116 349972 11172
rect 351148 16156 351204 16212
rect 352716 14364 352772 14420
rect 353612 6188 353668 6244
rect 354060 5852 354116 5908
rect 356188 17948 356244 18004
rect 359324 14588 359380 14644
rect 360332 16828 360388 16884
rect 357756 9212 357812 9268
rect 357868 9324 357924 9380
rect 354508 5852 354564 5908
rect 355964 6076 356020 6132
rect 364028 16828 364084 16884
rect 365372 16828 365428 16884
rect 362460 12572 362516 12628
rect 360892 11004 360948 11060
rect 360332 7980 360388 8036
rect 361676 7532 361732 7588
rect 359772 4396 359828 4452
rect 368732 17836 368788 17892
rect 367948 15932 368004 15988
rect 365596 9436 365652 9492
rect 367948 15708 368004 15764
rect 365372 2940 365428 2996
rect 365484 6300 365540 6356
rect 363580 2492 363636 2548
rect 367388 5964 367444 6020
rect 369628 5964 369684 6020
rect 371308 4284 371364 4340
rect 373436 16268 373492 16324
rect 374108 17724 374164 17780
rect 374108 14476 374164 14532
rect 371420 2604 371476 2660
rect 373100 14252 373156 14308
rect 376572 17724 376628 17780
rect 377132 17948 377188 18004
rect 375676 10892 375732 10948
rect 375004 10780 375060 10836
rect 376908 6188 376964 6244
rect 379708 16828 379764 16884
rect 378140 14252 378196 14308
rect 377132 6076 377188 6132
rect 378028 12684 378084 12740
rect 382844 17948 382900 18004
rect 379708 7644 379764 7700
rect 380716 7868 380772 7924
rect 385980 18060 386036 18116
rect 383516 16828 383572 16884
rect 383516 13020 383572 13076
rect 383068 7532 383124 7588
rect 384524 7756 384580 7812
rect 382620 4172 382676 4228
rect 387996 17612 388052 17668
rect 386428 2492 386484 2548
rect 386540 14364 386596 14420
rect 387996 14364 388052 14420
rect 388108 12796 388164 12852
rect 388892 17724 388948 17780
rect 388892 12908 388948 12964
rect 389788 14476 389844 14532
rect 388220 7868 388276 7924
rect 392252 16156 392308 16212
rect 390684 14476 390740 14532
rect 391468 16044 391524 16100
rect 393148 6300 393204 6356
rect 394044 11116 394100 11172
rect 395388 9324 395444 9380
rect 396508 14364 396564 14420
rect 395948 7980 396004 8036
rect 398524 17724 398580 17780
rect 400092 16044 400148 16100
rect 400652 17948 400708 18004
rect 396956 12796 397012 12852
rect 403228 17948 403284 18004
rect 401660 17612 401716 17668
rect 404796 14364 404852 14420
rect 404908 14588 404964 14644
rect 400652 6412 400708 6468
rect 403564 9212 403620 9268
rect 401660 6076 401716 6132
rect 399868 5852 399924 5908
rect 407932 18172 407988 18228
rect 407596 18060 407652 18116
rect 406364 9212 406420 9268
rect 407372 11004 407428 11060
rect 409500 12684 409556 12740
rect 407596 11004 407652 11060
rect 408268 12572 408324 12628
rect 412076 18172 412132 18228
rect 412636 11340 412692 11396
rect 412076 9548 412132 9604
rect 413084 9436 413140 9492
rect 409948 2716 410004 2772
rect 411180 2940 411236 2996
rect 413308 5852 413364 5908
rect 414092 17836 414148 17892
rect 415772 16828 415828 16884
rect 414092 5404 414148 5460
rect 414988 15932 415044 15988
rect 418348 15932 418404 15988
rect 418908 11228 418964 11284
rect 419132 16828 419188 16884
rect 420476 16828 420532 16884
rect 419132 6188 419188 6244
rect 421708 16268 421764 16324
rect 418796 5964 418852 6020
rect 416892 5404 416948 5460
rect 420700 2604 420756 2660
rect 422044 14700 422100 14756
rect 423612 12572 423668 12628
rect 424508 10892 424564 10948
rect 426748 17836 426804 17892
rect 427308 16828 427364 16884
rect 425180 12908 425236 12964
rect 427308 12908 427364 12964
rect 428428 14252 428484 14308
rect 426748 2604 426804 2660
rect 429884 14252 429940 14308
rect 430108 6076 430164 6132
rect 430220 13020 430276 13076
rect 433020 10892 433076 10948
rect 436156 16828 436212 16884
rect 433468 7756 433524 7812
rect 432124 7644 432180 7700
rect 435932 7532 435988 7588
rect 434028 6412 434084 6468
rect 439292 18172 439348 18228
rect 440860 16380 440916 16436
rect 440972 16828 441028 16884
rect 436828 7532 436884 7588
rect 437836 11004 437892 11060
rect 440972 7868 441028 7924
rect 441644 7980 441700 8036
rect 439740 2492 439796 2548
rect 443996 18060 444052 18116
rect 444332 17948 444388 18004
rect 441868 2492 441924 2548
rect 443548 14476 443604 14532
rect 444332 7980 444388 8036
rect 445228 16156 445284 16212
rect 445340 7644 445396 7700
rect 448700 17948 448756 18004
rect 449372 17724 449428 17780
rect 449260 9324 449316 9380
rect 447356 6300 447412 6356
rect 448812 5906 448868 5908
rect 448812 5854 448814 5906
rect 448814 5854 448866 5906
rect 448866 5854 448868 5906
rect 448812 5852 448868 5854
rect 450268 17724 450324 17780
rect 450380 18172 450436 18228
rect 453404 18172 453460 18228
rect 454972 16268 455028 16324
rect 456092 17612 456148 17668
rect 451836 14476 451892 14532
rect 453628 16044 453684 16100
rect 450380 13020 450436 13076
rect 449372 5068 449428 5124
rect 450268 12796 450324 12852
rect 425404 28 425460 84
rect 453068 5068 453124 5124
rect 458108 17612 458164 17668
rect 459228 17948 459284 18004
rect 456540 16156 456596 16212
rect 459676 14588 459732 14644
rect 459228 9436 459284 9492
rect 460348 14364 460404 14420
rect 458780 7980 458836 8036
rect 456092 6636 456148 6692
rect 456988 6636 457044 6692
rect 456204 6018 456260 6020
rect 456204 5966 456206 6018
rect 456206 5966 456258 6018
rect 456258 5966 456260 6018
rect 456204 5964 456260 5966
rect 456316 5906 456372 5908
rect 456316 5854 456318 5906
rect 456318 5854 456370 5906
rect 456370 5854 456372 5906
rect 456316 5852 456372 5854
rect 461244 11004 461300 11060
rect 464380 17948 464436 18004
rect 464604 18172 464660 18228
rect 464492 9548 464548 9604
rect 462028 4732 462084 4788
rect 462588 9212 462644 9268
rect 464604 2828 464660 2884
rect 465388 12684 465444 12740
rect 465948 11116 466004 11172
rect 467852 18060 467908 18116
rect 470652 18508 470708 18564
rect 469084 12796 469140 12852
rect 467852 6300 467908 6356
rect 470204 11340 470260 11396
rect 467068 4844 467124 4900
rect 468300 2716 468356 2772
rect 472108 5852 472164 5908
rect 475356 18060 475412 18116
rect 473788 16828 473844 16884
rect 475468 15932 475524 15988
rect 472220 4620 472276 4676
rect 474012 6188 474068 6244
rect 477932 17836 477988 17892
rect 475580 4508 475636 4564
rect 477820 11228 477876 11284
rect 478492 14364 478548 14420
rect 477932 6188 477988 6244
rect 478828 12908 478884 12964
rect 481628 17836 481684 17892
rect 480844 16828 480900 16884
rect 480060 9212 480116 9268
rect 480508 14700 480564 14756
rect 483196 12684 483252 12740
rect 484652 18060 484708 18116
rect 480844 9324 480900 9380
rect 482188 12572 482244 12628
rect 484764 12572 484820 12628
rect 489468 16828 489524 16884
rect 487228 5852 487284 5908
rect 487340 6188 487396 6244
rect 485548 4396 485604 4452
rect 484652 2716 484708 2772
rect 492604 18284 492660 18340
rect 492156 16828 492212 16884
rect 492156 16044 492212 16100
rect 490588 4284 490644 4340
rect 490700 14252 490756 14308
rect 489244 2604 489300 2660
rect 485772 28 485828 84
rect 495740 18060 495796 18116
rect 496412 17836 496468 17892
rect 494172 10780 494228 10836
rect 494956 10892 495012 10948
rect 493052 6076 493108 6132
rect 498876 18172 498932 18228
rect 497308 15932 497364 15988
rect 498092 17612 498148 17668
rect 496412 7756 496468 7812
rect 496860 7868 496916 7924
rect 498092 7868 498148 7924
rect 498764 7980 498820 8036
rect 502012 17836 502068 17892
rect 503132 17948 503188 18004
rect 501452 17724 501508 17780
rect 498988 4172 499044 4228
rect 500668 7532 500724 7588
rect 501452 6188 501508 6244
rect 502572 13020 502628 13076
rect 523292 532924 523348 532980
rect 521612 362908 521668 362964
rect 523292 430108 523348 430164
rect 556892 540988 556948 541044
rect 545132 536172 545188 536228
rect 540092 534380 540148 534436
rect 535052 531244 535108 531300
rect 533372 526092 533428 526148
rect 526652 112588 526708 112644
rect 530908 522732 530964 522788
rect 522508 20076 522564 20132
rect 519372 19964 519428 20020
rect 505148 17612 505204 17668
rect 506492 18284 506548 18340
rect 504028 14252 504084 14308
rect 504140 16380 504196 16436
rect 503132 6076 503188 6132
rect 513212 18172 513268 18228
rect 506492 7532 506548 7588
rect 510188 7644 510244 7700
rect 508284 6300 508340 6356
rect 506380 2492 506436 2548
rect 512092 5964 512148 6020
rect 520828 16268 520884 16324
rect 517468 14476 517524 14532
rect 513212 5964 513268 6020
rect 514108 9436 514164 9492
rect 515900 6188 515956 6244
rect 519708 2828 519764 2884
rect 522508 16156 522564 16212
rect 525868 14588 525924 14644
rect 525420 7868 525476 7924
rect 529228 11004 529284 11060
rect 538412 530908 538468 530964
rect 536732 529676 536788 529732
rect 536732 509068 536788 509124
rect 535052 468748 535108 468804
rect 533372 270508 533428 270564
rect 541772 519372 541828 519428
rect 553532 535948 553588 536004
rect 548492 532812 548548 532868
rect 550172 524524 550228 524580
rect 551852 521164 551908 521220
rect 551852 495628 551908 495684
rect 550172 416668 550228 416724
rect 548492 389788 548548 389844
rect 545132 349468 545188 349524
rect 541772 231868 541828 231924
rect 540092 191548 540148 191604
rect 538412 151228 538468 151284
rect 555212 525868 555268 525924
rect 560252 539532 560308 539588
rect 556892 310828 556948 310884
rect 558572 539420 558628 539476
rect 563612 536060 563668 536116
rect 566972 529452 567028 529508
rect 566972 455308 567028 455364
rect 563612 336028 563668 336084
rect 560252 297388 560308 297444
rect 558572 257068 558628 257124
rect 570332 551180 570388 551236
rect 580412 539308 580468 539364
rect 575372 537852 575428 537908
rect 575372 376348 575428 376404
rect 590492 527996 590548 528052
rect 589596 524412 589652 524468
rect 589596 522732 589652 522788
rect 593068 552748 593124 552804
rect 590604 523404 590660 523460
rect 590828 548940 590884 548996
rect 590828 523292 590884 523348
rect 590492 324492 590548 324548
rect 580412 218540 580468 218596
rect 570332 178108 570388 178164
rect 568652 137788 568708 137844
rect 555212 99148 555268 99204
rect 553532 58828 553588 58884
rect 593516 551068 593572 551124
rect 593404 546028 593460 546084
rect 593180 542780 593236 542836
rect 593180 483084 593236 483140
rect 593292 529228 593348 529284
rect 593068 33740 593124 33796
rect 593852 549388 593908 549444
rect 593628 524188 593684 524244
rect 593740 520828 593796 520884
rect 594412 541212 594468 541268
rect 594188 527548 594244 527604
rect 593964 520940 594020 520996
rect 594076 519260 594132 519316
rect 594300 525980 594356 526036
rect 594412 443436 594468 443492
rect 594524 519148 594580 519204
rect 594300 403788 594356 403844
rect 594188 284844 594244 284900
rect 594076 245196 594132 245252
rect 593964 205548 594020 205604
rect 593852 165900 593908 165956
rect 593740 126252 593796 126308
rect 593628 86604 593684 86660
rect 593516 73388 593572 73444
rect 593404 46956 593460 47012
rect 593292 20524 593348 20580
rect 539308 18508 539364 18564
rect 531468 18060 531524 18116
rect 537628 12796 537684 12852
rect 531468 11004 531524 11060
rect 534940 11116 534996 11172
rect 530908 8428 530964 8484
rect 533036 6076 533092 6132
rect 531132 4732 531188 4788
rect 536844 4844 536900 4900
rect 548492 17836 548548 17892
rect 544460 9324 544516 9380
rect 542668 4620 542724 4676
rect 577052 17612 577108 17668
rect 562828 16044 562884 16100
rect 548492 7644 548548 7700
rect 549388 14364 549444 14420
rect 548268 4508 548324 4564
rect 546364 2716 546420 2772
rect 554428 12684 554484 12740
rect 552076 9212 552132 9268
rect 553980 7756 554036 7812
rect 557788 12572 557844 12628
rect 561036 5852 561092 5908
rect 559692 4396 559748 4452
rect 573020 15932 573076 15988
rect 571228 11004 571284 11060
rect 569212 10892 569268 10948
rect 567308 7532 567364 7588
rect 565404 4284 565460 4340
rect 574924 5964 574980 6020
rect 581308 14252 581364 14308
rect 577052 4732 577108 4788
rect 580636 7644 580692 7700
rect 576828 4172 576884 4228
rect 594524 7308 594580 7364
rect 584444 4732 584500 4788
<< metal3 >>
rect 242722 593292 242732 593348
rect 242788 593292 496412 593348
rect 496468 593292 496478 593348
rect 234322 593180 234332 593236
rect 234388 593180 518476 593236
rect 518532 593180 518542 593236
rect 220882 593068 220892 593124
rect 220948 593068 584668 593124
rect 584724 593068 584734 593124
rect 335122 590604 335132 590660
rect 335188 590604 364028 590660
rect 364084 590604 364094 590660
rect 365362 590604 365372 590660
rect 365428 590604 452284 590660
rect 452340 590604 452350 590660
rect 261202 590492 261212 590548
rect 261268 590492 386092 590548
rect 386148 590492 386158 590548
rect 496402 590492 496412 590548
rect 496468 590492 562604 590548
rect 562660 590492 562670 590548
rect 165666 590156 165676 590212
rect 165732 590156 167132 590212
rect 167188 590156 167198 590212
rect 187730 590156 187740 590212
rect 187796 590156 188972 590212
rect 189028 590156 189038 590212
rect 253922 588812 253932 588868
rect 253988 588812 283948 588868
rect 284004 588812 284014 588868
rect 595560 588644 597000 588840
rect 590594 588588 590604 588644
rect 590660 588616 597000 588644
rect 590660 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 532 587188
rect 392 587132 532 587160
rect 476 587076 532 587132
rect 364 587020 532 587076
rect 364 586404 420 587020
rect 364 586348 337708 586404
rect 337764 586348 337774 586404
rect 274642 578732 274652 578788
rect 274708 578732 319228 578788
rect 319284 578732 319294 578788
rect 31938 577052 31948 577108
rect 32004 577052 332668 577108
rect 332724 577052 332734 577108
rect 595560 575428 597000 575624
rect 595420 575400 597000 575428
rect 595420 575372 595672 575400
rect 595420 575316 595476 575372
rect 595420 575260 595700 575316
rect 595644 574644 595700 575260
rect 232642 574588 232652 574644
rect 232708 574588 595700 574644
rect -960 573076 480 573272
rect -960 573048 8428 573076
rect 392 573020 8428 573048
rect 8372 572964 8428 573020
rect 8372 572908 346108 572964
rect 346164 572908 346174 572964
rect 280578 572012 280588 572068
rect 280644 572012 297388 572068
rect 297444 572012 297454 572068
rect 99138 570332 99148 570388
rect 99204 570332 319228 570388
rect 319284 570332 319294 570388
rect 167122 568652 167132 568708
rect 167188 568652 305788 568708
rect 305844 568652 305854 568708
rect 188962 566972 188972 567028
rect 189028 566972 297388 567028
rect 297444 566972 297454 567028
rect 267138 565292 267148 565348
rect 267204 565292 335132 565348
rect 335188 565292 335198 565348
rect 253698 563612 253708 563668
rect 253764 563612 430108 563668
rect 430164 563612 430174 563668
rect 595560 562212 597000 562408
rect 595420 562184 597000 562212
rect 595420 562156 595672 562184
rect 595420 562100 595476 562156
rect 595420 562044 595700 562100
rect 262098 561932 262108 561988
rect 262164 561932 341068 561988
rect 341124 561932 341134 561988
rect 595644 561204 595700 562044
rect 343522 561148 343532 561204
rect 343588 561148 595700 561204
rect 53778 560252 53788 560308
rect 53844 560252 324268 560308
rect 324324 560252 324334 560308
rect -960 558964 480 559160
rect -960 558936 532 558964
rect 392 558908 532 558936
rect 476 558852 532 558908
rect 364 558796 532 558852
rect 364 557844 420 558796
rect 364 557788 341068 557844
rect 341124 557788 341134 557844
rect 10098 556892 10108 556948
rect 10164 556892 327628 556948
rect 327684 556892 327694 556948
rect 5842 556108 5852 556164
rect 5908 556108 490588 556164
rect 490644 556108 490654 556164
rect 223458 555212 223468 555268
rect 223524 555212 539308 555268
rect 539364 555212 539374 555268
rect 17714 554428 17724 554484
rect 17780 554428 450268 554484
rect 450324 554428 450334 554484
rect 245298 553532 245308 553588
rect 245364 553532 365372 553588
rect 365428 553532 365438 553588
rect 70578 552860 70588 552916
rect 70644 552860 568652 552916
rect 568708 552860 568718 552916
rect 26898 552748 26908 552804
rect 26964 552748 593068 552804
rect 593124 552748 593134 552804
rect 228498 551852 228508 551908
rect 228564 551852 496412 551908
rect 496468 551852 496478 551908
rect 84018 551180 84028 551236
rect 84084 551180 570332 551236
rect 570388 551180 570398 551236
rect 40338 551068 40348 551124
rect 40404 551068 593516 551124
rect 593572 551068 593582 551124
rect 77298 550172 77308 550228
rect 77364 550172 315868 550228
rect 315924 550172 315934 550228
rect 19282 549500 19292 549556
rect 19348 549500 477148 549556
rect 477204 549500 477214 549556
rect 75618 549388 75628 549444
rect 75684 549388 593852 549444
rect 593908 549388 593918 549444
rect 595560 548996 597000 549192
rect 590818 548940 590828 548996
rect 590884 548968 597000 548996
rect 590884 548940 595672 548968
rect 206658 548492 206668 548548
rect 206724 548492 343532 548548
rect 343588 548492 343598 548548
rect 12562 547820 12572 547876
rect 12628 547820 480508 547876
rect 480564 547820 480574 547876
rect 2482 547708 2492 547764
rect 2548 547708 498988 547764
rect 499044 547708 499054 547764
rect 142818 546812 142828 546868
rect 142884 546812 302428 546868
rect 302484 546812 302494 546868
rect 15922 546140 15932 546196
rect 15988 546140 472108 546196
rect 472164 546140 472174 546196
rect 35298 546028 35308 546084
rect 35364 546028 593404 546084
rect 593460 546028 593470 546084
rect -960 544852 480 545048
rect -960 544824 532 544852
rect 392 544796 532 544824
rect 476 544740 532 544796
rect 364 544684 532 544740
rect 364 544516 420 544684
rect 19394 544572 19404 544628
rect 19460 544572 468748 544628
rect 468804 544572 468814 544628
rect 364 544460 349468 544516
rect 349524 544460 349534 544516
rect 53778 544348 53788 544404
rect 53844 544348 526652 544404
rect 526708 544348 526718 544404
rect 208338 543452 208348 543508
rect 208404 543452 288988 543508
rect 289044 543452 289054 543508
rect 9426 542892 9436 542948
rect 9492 542892 414988 542948
rect 415044 542892 415054 542948
rect 179778 542780 179788 542836
rect 179844 542780 593180 542836
rect 593236 542780 593246 542836
rect 9202 542668 9212 542724
rect 9268 542668 485548 542724
rect 485604 542668 485614 542724
rect 215058 541772 215068 541828
rect 215124 541772 232652 541828
rect 232708 541772 232718 541828
rect 250338 541772 250348 541828
rect 250404 541772 408268 541828
rect 408324 541772 408334 541828
rect 166338 541212 166348 541268
rect 166404 541212 594412 541268
rect 594468 541212 594478 541268
rect 10882 541100 10892 541156
rect 10948 541100 441868 541156
rect 441924 541100 441934 541156
rect 119298 540988 119308 541044
rect 119364 540988 556892 541044
rect 556948 540988 556958 541044
rect 14466 539644 14476 539700
rect 14532 539644 411628 539700
rect 411684 539644 411694 539700
rect 122658 539532 122668 539588
rect 122724 539532 560252 539588
rect 560308 539532 560318 539588
rect 109218 539420 109228 539476
rect 109284 539420 558572 539476
rect 558628 539420 558638 539476
rect 97458 539308 97468 539364
rect 97524 539308 580412 539364
rect 580468 539308 580478 539364
rect 17826 537964 17836 538020
rect 17892 537964 425068 538020
rect 425124 537964 425134 538020
rect 149538 537852 149548 537908
rect 149604 537852 575372 537908
rect 575428 537852 575438 537908
rect 10994 537740 11004 537796
rect 11060 537740 436828 537796
rect 436884 537740 436894 537796
rect 5954 537628 5964 537684
rect 6020 537628 463708 537684
rect 463764 537628 463774 537684
rect 14690 536284 14700 536340
rect 14756 536284 371868 536340
rect 371924 536284 371934 536340
rect 131618 536172 131628 536228
rect 131684 536172 545132 536228
rect 545188 536172 545198 536228
rect 136098 536060 136108 536116
rect 136164 536060 563612 536116
rect 563668 536060 563678 536116
rect 44258 535948 44268 536004
rect 44324 535948 553532 536004
rect 553588 535948 553598 536004
rect 595560 535780 597000 535976
rect 595420 535752 597000 535780
rect 595420 535724 595672 535752
rect 595420 535668 595476 535724
rect 595420 535612 595700 535668
rect 141250 534604 141260 534660
rect 141316 534604 521612 534660
rect 521668 534604 521678 534660
rect 2706 534492 2716 534548
rect 2772 534492 398188 534548
rect 398244 534492 398254 534548
rect 79202 534380 79212 534436
rect 79268 534380 540092 534436
rect 540148 534380 540158 534436
rect 595644 534324 595700 535612
rect 201618 534268 201628 534324
rect 201684 534268 595700 534324
rect 157938 532924 157948 532980
rect 158004 532924 523292 532980
rect 523348 532924 523358 532980
rect 144722 532812 144732 532868
rect 144788 532812 548492 532868
rect 548548 532812 548558 532868
rect 14354 532700 14364 532756
rect 14420 532700 459228 532756
rect 459284 532700 459294 532756
rect 130 532588 140 532644
rect 196 532588 447020 532644
rect 447076 532588 447086 532644
rect 171378 531244 171388 531300
rect 171444 531244 535052 531300
rect 535108 531244 535118 531300
rect 11106 531132 11116 531188
rect 11172 531132 393708 531188
rect 393764 531132 393774 531188
rect 17602 531020 17612 531076
rect 17668 531020 455308 531076
rect 455364 531020 455374 531076
rect -960 530740 480 530936
rect 66098 530908 66108 530964
rect 66164 530908 538412 530964
rect 538468 530908 538478 530964
rect -960 530712 532 530740
rect 392 530684 532 530712
rect 476 530628 532 530684
rect 364 530572 532 530628
rect 364 529396 420 530572
rect 184930 529676 184940 529732
rect 184996 529676 536732 529732
rect 536788 529676 536798 529732
rect 9314 529564 9324 529620
rect 9380 529564 389788 529620
rect 389844 529564 389854 529620
rect 175298 529452 175308 529508
rect 175364 529452 566972 529508
rect 567028 529452 567038 529508
rect 364 529340 359660 529396
rect 359716 529340 359726 529396
rect 32050 529228 32060 529284
rect 32116 529228 593292 529284
rect 593348 529228 593358 529284
rect 231858 527996 231868 528052
rect 231924 527996 590492 528052
rect 590548 527996 590558 528052
rect 12786 527884 12796 527940
rect 12852 527884 385084 527940
rect 385140 527884 385150 527940
rect 19506 527772 19516 527828
rect 19572 527772 403340 527828
rect 403396 527772 403406 527828
rect 2594 527660 2604 527716
rect 2660 527660 420028 527716
rect 420084 527660 420094 527716
rect 115602 527548 115612 527604
rect 115668 527548 594188 527604
rect 594244 527548 594254 527604
rect 16146 526316 16156 526372
rect 16212 526316 381500 526372
rect 381556 526316 381566 526372
rect 12674 526204 12684 526260
rect 12740 526204 406924 526260
rect 406980 526204 406990 526260
rect 106866 526092 106876 526148
rect 106932 526092 533372 526148
rect 533428 526092 533438 526148
rect 154466 525980 154476 526036
rect 154532 525980 594300 526036
rect 594356 525980 594366 526036
rect 58482 525868 58492 525924
rect 58548 525868 555212 525924
rect 555268 525868 555278 525924
rect 5058 524636 5068 524692
rect 5124 524636 354508 524692
rect 354564 524636 354574 524692
rect 163650 524524 163660 524580
rect 163716 524524 550172 524580
rect 550228 524524 550238 524580
rect 194226 524412 194236 524468
rect 194292 524412 589596 524468
rect 589652 524412 589662 524468
rect 16034 524300 16044 524356
rect 16100 524300 428764 524356
rect 428820 524300 428830 524356
rect 50082 524188 50092 524244
rect 50148 524188 593628 524244
rect 593684 524188 593694 524244
rect 230178 523740 230188 523796
rect 230244 523740 294140 523796
rect 294196 523740 294206 523796
rect 120978 523628 120988 523684
rect 121044 523628 310828 523684
rect 310884 523628 310894 523684
rect 128706 523516 128716 523572
rect 128772 523516 231868 523572
rect 231924 523516 231934 523572
rect 237906 523516 237916 523572
rect 237972 523516 473788 523572
rect 473844 523516 473854 523572
rect 211586 523404 211596 523460
rect 211652 523404 590604 523460
rect 590660 523404 590670 523460
rect 198146 523292 198156 523348
rect 198212 523292 590828 523348
rect 590884 523292 590894 523348
rect 219874 523180 219884 523236
rect 219940 523180 220892 523236
rect 220948 523180 220958 523236
rect 233426 522732 233436 522788
rect 233492 522732 234332 522788
rect 234388 522732 234398 522788
rect 241826 522732 241836 522788
rect 241892 522732 242732 522788
rect 242788 522732 242798 522788
rect 259746 522732 259756 522788
rect 259812 522732 261212 522788
rect 261268 522732 261278 522788
rect 272738 522732 272748 522788
rect 272804 522732 274652 522788
rect 274708 522732 274718 522788
rect 513090 522732 513100 522788
rect 513156 522732 530908 522788
rect 530964 522732 530974 522788
rect 589586 522732 589596 522788
rect 589652 522760 595672 522788
rect 589652 522732 597000 522760
rect 14578 522620 14588 522676
rect 14644 522620 367948 522676
rect 368004 522620 368014 522676
rect 508722 522620 508732 522676
rect 508788 522620 519372 522676
rect 519428 522620 519438 522676
rect 14242 522508 14252 522564
rect 14308 522508 503020 522564
rect 503076 522508 503086 522564
rect 595560 522536 597000 522732
rect 9538 521276 9548 521332
rect 9604 521276 363244 521332
rect 363300 521276 363310 521332
rect 189746 521164 189756 521220
rect 189812 521164 551852 521220
rect 551908 521164 551918 521220
rect 18 521052 28 521108
rect 84 521052 494284 521108
rect 494340 521052 494350 521108
rect 88946 520940 88956 520996
rect 89012 520940 593964 520996
rect 594020 520940 594030 520996
rect 63186 520828 63196 520884
rect 63252 520828 593740 520884
rect 593796 520828 593806 520884
rect 19618 519596 19628 519652
rect 19684 519596 377020 519652
rect 377076 519596 377086 519652
rect 6066 519484 6076 519540
rect 6132 519484 433804 519540
rect 433860 519484 433870 519540
rect 93090 519372 93100 519428
rect 93156 519372 541772 519428
rect 541828 519372 541838 519428
rect 23202 519260 23212 519316
rect 23268 519260 31948 519316
rect 101826 519260 101836 519316
rect 101892 519260 594076 519316
rect 594132 519260 594142 519316
rect 31892 519204 31948 519260
rect 31892 519148 594524 519204
rect 594580 519148 594590 519204
rect 392 516824 5068 516852
rect -960 516796 5068 516824
rect 5124 516796 5134 516852
rect -960 516600 480 516796
rect 595560 509348 597000 509544
rect 572852 509320 597000 509348
rect 572852 509292 595672 509320
rect 572852 509124 572908 509292
rect 536722 509068 536732 509124
rect 536788 509068 572908 509124
rect 392 502712 9548 502740
rect -960 502684 9548 502712
rect 9604 502684 9614 502740
rect -960 502488 480 502684
rect 595560 496132 597000 496328
rect 595420 496104 597000 496132
rect 595420 496076 595672 496104
rect 595420 496020 595476 496076
rect 595420 495964 595700 496020
rect 595644 495684 595700 495964
rect 551842 495628 551852 495684
rect 551908 495628 595700 495684
rect -960 488404 480 488600
rect -960 488376 532 488404
rect 392 488348 532 488376
rect 476 488292 532 488348
rect 364 488236 532 488292
rect 364 487284 420 488236
rect 364 487228 14700 487284
rect 14756 487228 14766 487284
rect 593170 483084 593180 483140
rect 593236 483112 595672 483140
rect 593236 483084 597000 483112
rect 595560 482888 597000 483084
rect -960 474292 480 474488
rect -960 474264 532 474292
rect 392 474236 532 474264
rect 476 474180 532 474236
rect 364 474124 532 474180
rect 364 473844 420 474124
rect 364 473788 14588 473844
rect 14644 473788 14654 473844
rect 595560 469700 597000 469896
rect 595420 469672 597000 469700
rect 595420 469644 595672 469672
rect 595420 469588 595476 469644
rect 595420 469532 595700 469588
rect 595644 468804 595700 469532
rect 535042 468748 535052 468804
rect 535108 468748 595700 468804
rect -960 460180 480 460376
rect -960 460152 532 460180
rect 392 460124 532 460152
rect 476 460068 532 460124
rect 364 460012 532 460068
rect 364 458724 420 460012
rect 364 458668 19628 458724
rect 19684 458668 19694 458724
rect 595560 456484 597000 456680
rect 595420 456456 597000 456484
rect 595420 456428 595672 456456
rect 595420 456372 595476 456428
rect 595420 456316 595700 456372
rect 595644 455364 595700 456316
rect 566962 455308 566972 455364
rect 567028 455308 595700 455364
rect -960 446068 480 446264
rect -960 446040 532 446068
rect 392 446012 532 446040
rect 476 445956 532 446012
rect 364 445900 532 445956
rect 364 445284 420 445900
rect 364 445228 12796 445284
rect 12852 445228 12862 445284
rect 594402 443436 594412 443492
rect 594468 443464 595672 443492
rect 594468 443436 597000 443464
rect 595560 443240 597000 443436
rect -960 431956 480 432152
rect -960 431928 16156 431956
rect 392 431900 16156 431928
rect 16212 431900 16222 431956
rect 595560 430164 597000 430248
rect 523282 430108 523292 430164
rect 523348 430108 597000 430164
rect 595560 430024 597000 430108
rect 392 418040 9324 418068
rect -960 418012 9324 418040
rect 9380 418012 9390 418068
rect -960 417816 480 418012
rect 595560 416836 597000 417032
rect 572852 416808 597000 416836
rect 572852 416780 595672 416808
rect 572852 416724 572908 416780
rect 550162 416668 550172 416724
rect 550228 416668 572908 416724
rect 392 403928 2716 403956
rect -960 403900 2716 403928
rect 2772 403900 2782 403956
rect -960 403704 480 403900
rect 594290 403788 594300 403844
rect 594356 403816 595672 403844
rect 594356 403788 597000 403816
rect 595560 403592 597000 403788
rect 595560 390404 597000 390600
rect 595420 390376 597000 390404
rect 595420 390348 595672 390376
rect 595420 390292 595476 390348
rect 595420 390236 595700 390292
rect 595644 389844 595700 390236
rect -960 389732 480 389816
rect 548482 389788 548492 389844
rect 548548 389788 595700 389844
rect -960 389676 11116 389732
rect 11172 389676 11182 389732
rect -960 389592 480 389676
rect 595560 377188 597000 377384
rect 595420 377160 597000 377188
rect 595420 377132 595672 377160
rect 595420 377076 595476 377132
rect 595420 377020 595700 377076
rect 595644 376404 595700 377020
rect 575362 376348 575372 376404
rect 575428 376348 595700 376404
rect -960 375508 480 375704
rect -960 375480 532 375508
rect 392 375452 532 375480
rect 476 375396 532 375452
rect 364 375340 532 375396
rect 364 374724 420 375340
rect 364 374668 19516 374724
rect 19572 374668 19582 374724
rect 595560 363972 597000 364168
rect 595420 363944 597000 363972
rect 595420 363916 595672 363944
rect 595420 363860 595476 363916
rect 595420 363804 595700 363860
rect 595644 362964 595700 363804
rect 521602 362908 521612 362964
rect 521668 362908 595700 362964
rect -960 361396 480 361592
rect -960 361368 14476 361396
rect 392 361340 14476 361368
rect 14532 361340 14542 361396
rect 595560 350756 597000 350952
rect 595420 350728 597000 350756
rect 595420 350700 595672 350728
rect 595420 350644 595476 350700
rect 595420 350588 595700 350644
rect 595644 349524 595700 350588
rect 545122 349468 545132 349524
rect 545188 349468 595700 349524
rect -960 347284 480 347480
rect -960 347256 532 347284
rect 392 347228 532 347256
rect 476 347172 532 347228
rect 364 347116 532 347172
rect 364 346164 420 347116
rect 364 346108 12684 346164
rect 12740 346108 12750 346164
rect 595560 337540 597000 337736
rect 595420 337512 597000 337540
rect 595420 337484 595672 337512
rect 595420 337428 595476 337484
rect 595420 337372 595700 337428
rect 595644 336084 595700 337372
rect 563602 336028 563612 336084
rect 563668 336028 595700 336084
rect 392 333368 9436 333396
rect -960 333340 9436 333368
rect 9492 333340 9502 333396
rect -960 333144 480 333340
rect 590482 324492 590492 324548
rect 590548 324520 595672 324548
rect 590548 324492 597000 324520
rect 595560 324296 597000 324492
rect -960 319060 480 319256
rect -960 319032 532 319060
rect 392 319004 532 319032
rect 476 318948 532 319004
rect 364 318892 532 318948
rect 364 317604 420 318892
rect 364 317548 17836 317604
rect 17892 317548 17902 317604
rect 595560 311108 597000 311304
rect 572852 311080 597000 311108
rect 572852 311052 595672 311080
rect 572852 310884 572908 311052
rect 556882 310828 556892 310884
rect 556948 310828 572908 310884
rect 392 305144 2604 305172
rect -960 305116 2604 305144
rect 2660 305116 2670 305172
rect -960 304920 480 305116
rect 595560 297892 597000 298088
rect 595420 297864 597000 297892
rect 595420 297836 595672 297864
rect 595420 297780 595476 297836
rect 595420 297724 595700 297780
rect 595644 297444 595700 297724
rect 560242 297388 560252 297444
rect 560308 297388 595700 297444
rect -960 290836 480 291032
rect -960 290808 16044 290836
rect 392 290780 16044 290808
rect 16100 290780 16110 290836
rect 594178 284844 594188 284900
rect 594244 284872 595672 284900
rect 594244 284844 597000 284872
rect 595560 284648 597000 284844
rect 392 276920 11004 276948
rect -960 276892 11004 276920
rect 11060 276892 11070 276948
rect -960 276696 480 276892
rect 595560 271460 597000 271656
rect 595420 271432 597000 271460
rect 595420 271404 595672 271432
rect 595420 271348 595476 271404
rect 595420 271292 595700 271348
rect 595644 270564 595700 271292
rect 533362 270508 533372 270564
rect 533428 270508 595700 270564
rect 392 262808 6076 262836
rect -960 262780 6076 262808
rect 6132 262780 6142 262836
rect -960 262584 480 262780
rect 595560 258244 597000 258440
rect 595420 258216 597000 258244
rect 595420 258188 595672 258216
rect 595420 258132 595476 258188
rect 595420 258076 595700 258132
rect 595644 257124 595700 258076
rect 558562 257068 558572 257124
rect 558628 257068 595700 257124
rect -960 248612 480 248696
rect -960 248556 10892 248612
rect 10948 248556 10958 248612
rect -960 248472 480 248556
rect 594066 245196 594076 245252
rect 594132 245224 595672 245252
rect 594132 245196 597000 245224
rect 595560 245000 597000 245196
rect -960 234388 480 234584
rect -960 234360 532 234388
rect 392 234332 532 234360
rect 476 234276 532 234332
rect 364 234220 532 234276
rect 364 233604 420 234220
rect 364 233548 17724 233604
rect 17780 233548 17790 233604
rect 595560 231924 597000 232008
rect 541762 231868 541772 231924
rect 541828 231868 597000 231924
rect 595560 231784 597000 231868
rect 130 220556 140 220612
rect 196 220556 532 220612
rect 476 220500 532 220556
rect 392 220472 532 220500
rect -960 220444 532 220472
rect -960 220248 480 220444
rect 595560 218596 597000 218792
rect 580402 218540 580412 218596
rect 580468 218568 597000 218596
rect 580468 218540 595672 218568
rect -960 206164 480 206360
rect -960 206136 532 206164
rect 392 206108 532 206136
rect 476 206052 532 206108
rect 364 205996 532 206052
rect 364 205044 420 205996
rect 593954 205548 593964 205604
rect 594020 205576 595672 205604
rect 594020 205548 597000 205576
rect 595560 205352 597000 205548
rect 364 204988 17612 205044
rect 17668 204988 17678 205044
rect 392 192248 5964 192276
rect -960 192220 5964 192248
rect 6020 192220 6030 192276
rect -960 192024 480 192220
rect 595560 192164 597000 192360
rect 595420 192136 597000 192164
rect 595420 192108 595672 192136
rect 595420 192052 595476 192108
rect 595420 191996 595700 192052
rect 595644 191604 595700 191996
rect 540082 191548 540092 191604
rect 540148 191548 595700 191604
rect 595560 178948 597000 179144
rect 595420 178920 597000 178948
rect 595420 178892 595672 178920
rect 595420 178836 595476 178892
rect 595420 178780 595700 178836
rect 595644 178164 595700 178780
rect -960 177940 480 178136
rect 570322 178108 570332 178164
rect 570388 178108 595700 178164
rect -960 177912 532 177940
rect 392 177884 532 177912
rect 476 177828 532 177884
rect 364 177772 532 177828
rect 364 176484 420 177772
rect 364 176428 14364 176484
rect 14420 176428 14430 176484
rect 593842 165900 593852 165956
rect 593908 165928 595672 165956
rect 593908 165900 597000 165928
rect 595560 165704 597000 165900
rect -960 163828 480 164024
rect -960 163800 532 163828
rect 392 163772 532 163800
rect 476 163716 532 163772
rect 364 163660 532 163716
rect 364 163044 420 163660
rect 364 162988 19404 163044
rect 19460 162988 19470 163044
rect 595560 152516 597000 152712
rect 595420 152488 597000 152516
rect 595420 152460 595672 152488
rect 595420 152404 595476 152460
rect 595420 152348 595700 152404
rect 595644 151284 595700 152348
rect 538402 151228 538412 151284
rect 538468 151228 595700 151284
rect -960 149716 480 149912
rect -960 149688 19292 149716
rect 392 149660 19292 149688
rect 19348 149660 19358 149716
rect 595560 139300 597000 139496
rect 595420 139272 597000 139300
rect 595420 139244 595672 139272
rect 595420 139188 595476 139244
rect 595420 139132 595700 139188
rect 595644 137844 595700 139132
rect 568642 137788 568652 137844
rect 568708 137788 595700 137844
rect -960 135604 480 135800
rect -960 135576 532 135604
rect 392 135548 532 135576
rect 476 135492 532 135548
rect 364 135436 532 135492
rect 364 134484 420 135436
rect 364 134428 15932 134484
rect 15988 134428 15998 134484
rect 593730 126252 593740 126308
rect 593796 126280 595672 126308
rect 593796 126252 597000 126280
rect 595560 126056 597000 126252
rect -960 121492 480 121688
rect -960 121464 532 121492
rect 392 121436 532 121464
rect 476 121380 532 121436
rect 364 121324 532 121380
rect 364 121044 420 121324
rect 364 120988 12572 121044
rect 12628 120988 12638 121044
rect 595560 112868 597000 113064
rect 572852 112840 597000 112868
rect 572852 112812 595672 112840
rect 572852 112644 572908 112812
rect 526642 112588 526652 112644
rect 526708 112588 572908 112644
rect -960 107492 480 107576
rect -960 107436 5852 107492
rect 5908 107436 5918 107492
rect -960 107352 480 107436
rect 595560 99652 597000 99848
rect 595420 99624 597000 99652
rect 595420 99596 595672 99624
rect 595420 99540 595476 99596
rect 595420 99484 595700 99540
rect 595644 99204 595700 99484
rect 555202 99148 555212 99204
rect 555268 99148 595700 99204
rect 392 93464 9212 93492
rect -960 93436 9212 93464
rect 9268 93436 9278 93492
rect -960 93240 480 93436
rect 593618 86604 593628 86660
rect 593684 86632 595672 86660
rect 593684 86604 597000 86632
rect 595560 86408 597000 86604
rect 18 79436 28 79492
rect 84 79436 532 79492
rect 476 79380 532 79436
rect 392 79352 532 79380
rect -960 79324 532 79352
rect -960 79128 480 79324
rect 593506 73388 593516 73444
rect 593572 73416 595672 73444
rect 593572 73388 597000 73416
rect 595560 73192 597000 73388
rect -960 65044 480 65240
rect -960 65016 532 65044
rect 392 64988 532 65016
rect 476 64932 532 64988
rect 364 64876 532 64932
rect 364 63924 420 64876
rect 364 63868 14252 63924
rect 14308 63868 14318 63924
rect 595560 60004 597000 60200
rect 595420 59976 597000 60004
rect 595420 59948 595672 59976
rect 595420 59892 595476 59948
rect 595420 59836 595700 59892
rect 595644 58884 595700 59836
rect 553522 58828 553532 58884
rect 553588 58828 595700 58884
rect 392 51128 2492 51156
rect -960 51100 2492 51128
rect 2548 51100 2558 51156
rect -960 50904 480 51100
rect 593394 46956 593404 47012
rect 593460 46984 595672 47012
rect 593460 46956 597000 46984
rect 595560 46760 597000 46956
rect -960 36820 480 37016
rect -960 36792 4172 36820
rect 392 36764 4172 36792
rect 4228 36764 4238 36820
rect 593058 33740 593068 33796
rect 593124 33768 595672 33796
rect 593124 33740 597000 33768
rect 595560 33544 597000 33740
rect -960 22708 480 22904
rect -960 22680 4956 22708
rect 392 22652 4956 22680
rect 5012 22652 5022 22708
rect 593282 20524 593292 20580
rect 593348 20552 595672 20580
rect 593348 20524 597000 20552
rect 595560 20328 597000 20524
rect 4946 20076 4956 20132
rect 5012 20076 522508 20132
rect 522564 20076 522574 20132
rect 4162 19964 4172 20020
rect 4228 19964 519372 20020
rect 519428 19964 519438 20020
rect 470642 18508 470652 18564
rect 470708 18508 539308 18564
rect 539364 18508 539374 18564
rect 97682 18396 97692 18452
rect 97748 18396 106204 18452
rect 106260 18396 106270 18452
rect 32722 18284 32732 18340
rect 32788 18284 43932 18340
rect 43988 18284 43998 18340
rect 92530 18284 92540 18340
rect 92596 18284 101500 18340
rect 101556 18284 101566 18340
rect 492594 18284 492604 18340
rect 492660 18284 506492 18340
rect 506548 18284 506558 18340
rect 40450 18172 40460 18228
rect 40516 18172 59164 18228
rect 59220 18172 59230 18228
rect 69010 18172 69020 18228
rect 69076 18172 82684 18228
rect 82740 18172 82750 18228
rect 90738 18172 90748 18228
rect 90804 18172 99932 18228
rect 99988 18172 99998 18228
rect 105858 18172 105868 18228
rect 105924 18172 112588 18228
rect 112644 18172 112654 18228
rect 407922 18172 407932 18228
rect 407988 18172 412076 18228
rect 412132 18172 412142 18228
rect 439282 18172 439292 18228
rect 439348 18172 450380 18228
rect 450436 18172 450446 18228
rect 453394 18172 453404 18228
rect 453460 18172 464604 18228
rect 464660 18172 464670 18228
rect 498866 18172 498876 18228
rect 498932 18172 513212 18228
rect 513268 18172 513278 18228
rect 33618 18060 33628 18116
rect 33684 18060 52892 18116
rect 52948 18060 52958 18116
rect 67218 18060 67228 18116
rect 67284 18060 81116 18116
rect 81172 18060 81182 18116
rect 102722 18060 102732 18116
rect 102788 18060 109340 18116
rect 109396 18060 109406 18116
rect 385970 18060 385980 18116
rect 386036 18060 407596 18116
rect 407652 18060 407662 18116
rect 443986 18060 443996 18116
rect 444052 18060 467852 18116
rect 467908 18060 467918 18116
rect 475346 18060 475356 18116
rect 475412 18060 484652 18116
rect 484708 18060 484718 18116
rect 495730 18060 495740 18116
rect 495796 18060 531468 18116
rect 531524 18060 531534 18116
rect 35298 17948 35308 18004
rect 35364 17948 54460 18004
rect 54516 17948 54526 18004
rect 63858 17948 63868 18004
rect 63924 17948 77980 18004
rect 78036 17948 78046 18004
rect 89058 17948 89068 18004
rect 89124 17948 98364 18004
rect 98420 17948 98430 18004
rect 104178 17948 104188 18004
rect 104244 17948 110908 18004
rect 110964 17948 110974 18004
rect 335794 17948 335804 18004
rect 335860 17948 353612 18004
rect 353668 17948 353678 18004
rect 356178 17948 356188 18004
rect 356244 17948 377132 18004
rect 377188 17948 377198 18004
rect 382834 17948 382844 18004
rect 382900 17948 400652 18004
rect 400708 17948 400718 18004
rect 403218 17948 403228 18004
rect 403284 17948 444332 18004
rect 444388 17948 444398 18004
rect 448690 17948 448700 18004
rect 448756 17948 459228 18004
rect 459284 17948 459294 18004
rect 464370 17948 464380 18004
rect 464436 17948 503132 18004
rect 503188 17948 503198 18004
rect 36978 17836 36988 17892
rect 37044 17836 56364 17892
rect 56420 17836 56430 17892
rect 62178 17836 62188 17892
rect 62244 17836 76412 17892
rect 76468 17836 76478 17892
rect 276210 17836 276220 17892
rect 276276 17836 289772 17892
rect 289828 17836 289838 17892
rect 291890 17836 291900 17892
rect 291956 17836 306908 17892
rect 306964 17836 306974 17892
rect 326386 17836 326396 17892
rect 326452 17836 346892 17892
rect 346948 17836 346958 17892
rect 368722 17836 368732 17892
rect 368788 17836 414092 17892
rect 414148 17836 414158 17892
rect 426738 17836 426748 17892
rect 426804 17836 477932 17892
rect 477988 17836 477998 17892
rect 481618 17836 481628 17892
rect 481684 17836 496412 17892
rect 496468 17836 496478 17892
rect 502002 17836 502012 17892
rect 502068 17836 548492 17892
rect 548548 17836 548558 17892
rect 38658 17724 38668 17780
rect 38724 17724 57596 17780
rect 57652 17724 57662 17780
rect 65538 17724 65548 17780
rect 65604 17724 79884 17780
rect 79940 17724 79950 17780
rect 85698 17724 85708 17780
rect 85764 17724 95788 17780
rect 95844 17724 95854 17780
rect 110898 17724 110908 17780
rect 110964 17724 117628 17780
rect 117684 17724 117694 17780
rect 290322 17724 290332 17780
rect 290388 17724 314972 17780
rect 315028 17724 315038 17780
rect 316978 17724 316988 17780
rect 317044 17724 343532 17780
rect 343588 17724 343598 17780
rect 346770 17724 346780 17780
rect 346836 17724 374108 17780
rect 374164 17724 374174 17780
rect 376562 17724 376572 17780
rect 376628 17724 388892 17780
rect 388948 17724 388958 17780
rect 398514 17724 398524 17780
rect 398580 17724 449372 17780
rect 449428 17724 449438 17780
rect 450258 17724 450268 17780
rect 450324 17724 501452 17780
rect 501508 17724 501518 17780
rect 18498 17612 18508 17668
rect 18564 17612 40348 17668
rect 40404 17612 40414 17668
rect 60498 17612 60508 17668
rect 60564 17612 74844 17668
rect 74900 17612 74910 17668
rect 87490 17612 87500 17668
rect 87556 17612 97468 17668
rect 97524 17612 97534 17668
rect 100818 17612 100828 17668
rect 100884 17612 107772 17668
rect 107828 17612 107838 17668
rect 114258 17612 114268 17668
rect 114324 17612 119308 17668
rect 119364 17612 119374 17668
rect 238578 17612 238588 17668
rect 238644 17612 257852 17668
rect 257908 17612 257918 17668
rect 260530 17612 260540 17668
rect 260596 17612 285516 17668
rect 285572 17612 285582 17668
rect 288754 17612 288764 17668
rect 288820 17612 308252 17668
rect 308308 17612 308318 17668
rect 309138 17612 309148 17668
rect 309204 17612 336812 17668
rect 336868 17612 336878 17668
rect 353042 17612 353052 17668
rect 353108 17612 387996 17668
rect 388052 17612 388062 17668
rect 401650 17612 401660 17668
rect 401716 17612 456092 17668
rect 456148 17612 456158 17668
rect 458098 17612 458108 17668
rect 458164 17612 498092 17668
rect 498148 17612 498158 17668
rect 505138 17612 505148 17668
rect 505204 17612 577052 17668
rect 577108 17612 577118 17668
rect 343634 17276 343644 17332
rect 343700 17276 352716 17332
rect 352772 17276 352782 17332
rect 273074 17164 273084 17220
rect 273140 17164 275436 17220
rect 275492 17164 275502 17220
rect 94098 16940 94108 16996
rect 94164 16940 103516 16996
rect 103572 16940 103582 16996
rect 107650 16940 107660 16996
rect 107716 16940 114492 16996
rect 114548 16940 114558 16996
rect 116050 16940 116060 16996
rect 116116 16940 120988 16996
rect 121044 16940 121054 16996
rect 95890 16828 95900 16884
rect 95956 16828 104636 16884
rect 104692 16828 104702 16884
rect 109218 16828 109228 16884
rect 109284 16828 115948 16884
rect 116004 16828 116014 16884
rect 257394 16828 257404 16884
rect 257460 16828 261212 16884
rect 261268 16828 261278 16884
rect 285618 16828 285628 16884
rect 285684 16828 288764 16884
rect 288820 16828 288830 16884
rect 295026 16828 295036 16884
rect 295092 16828 296492 16884
rect 296548 16828 296558 16884
rect 310706 16828 310716 16884
rect 310772 16828 312396 16884
rect 312452 16828 312462 16884
rect 313842 16828 313852 16884
rect 313908 16828 316652 16884
rect 316708 16828 316718 16884
rect 332658 16828 332668 16884
rect 332724 16828 335356 16884
rect 335412 16828 335422 16884
rect 351474 16828 351484 16884
rect 351540 16828 360332 16884
rect 360388 16828 360398 16884
rect 364018 16828 364028 16884
rect 364084 16828 365372 16884
rect 365428 16828 365438 16884
rect 379698 16828 379708 16884
rect 379764 16828 383516 16884
rect 383572 16828 383582 16884
rect 415762 16828 415772 16884
rect 415828 16828 419132 16884
rect 419188 16828 419198 16884
rect 420466 16828 420476 16884
rect 420532 16828 427308 16884
rect 427364 16828 427374 16884
rect 436146 16828 436156 16884
rect 436212 16828 440972 16884
rect 441028 16828 441038 16884
rect 473778 16828 473788 16884
rect 473844 16828 480844 16884
rect 480900 16828 480910 16884
rect 489458 16828 489468 16884
rect 489524 16828 492156 16884
rect 492212 16828 492222 16884
rect 216626 16492 216636 16548
rect 216692 16492 231868 16548
rect 231924 16492 231934 16548
rect 224466 16380 224476 16436
rect 224532 16380 240268 16436
rect 240324 16380 240334 16436
rect 440850 16380 440860 16436
rect 440916 16380 504140 16436
rect 504196 16380 504206 16436
rect 221330 16268 221340 16324
rect 221396 16268 236908 16324
rect 236964 16268 236974 16324
rect 373426 16268 373436 16324
rect 373492 16268 421708 16324
rect 421764 16268 421774 16324
rect 454962 16268 454972 16324
rect 455028 16268 520828 16324
rect 520884 16268 520894 16324
rect 222898 16156 222908 16212
rect 222964 16156 238588 16212
rect 238644 16156 238654 16212
rect 315410 16156 315420 16212
rect 315476 16156 351148 16212
rect 351204 16156 351214 16212
rect 392242 16156 392252 16212
rect 392308 16156 445228 16212
rect 445284 16156 445294 16212
rect 456530 16156 456540 16212
rect 456596 16156 522508 16212
rect 522564 16156 522574 16212
rect 218194 16044 218204 16100
rect 218260 16044 233548 16100
rect 233604 16044 233614 16100
rect 246418 16044 246428 16100
rect 246484 16044 267148 16100
rect 267204 16044 267214 16100
rect 271506 16044 271516 16100
rect 271572 16044 297388 16100
rect 297444 16044 297454 16100
rect 349458 16044 349468 16100
rect 349524 16044 391468 16100
rect 391524 16044 391534 16100
rect 400082 16044 400092 16100
rect 400148 16044 453628 16100
rect 453684 16044 453694 16100
rect 492146 16044 492156 16100
rect 492212 16044 562828 16100
rect 562884 16044 562894 16100
rect 30370 15932 30380 15988
rect 30436 15932 50428 15988
rect 50484 15932 50494 15988
rect 219762 15932 219772 15988
rect 219828 15932 235228 15988
rect 235284 15932 235294 15988
rect 262098 15932 262108 15988
rect 262164 15932 287420 15988
rect 287476 15932 287486 15988
rect 288754 15932 288764 15988
rect 288820 15932 315980 15988
rect 316036 15932 316046 15988
rect 329522 15932 329532 15988
rect 329588 15932 361228 15988
rect 367938 15932 367948 15988
rect 368004 15932 414988 15988
rect 415044 15932 415054 15988
rect 418338 15932 418348 15988
rect 418404 15932 475468 15988
rect 475524 15932 475534 15988
rect 497298 15932 497308 15988
rect 497364 15932 573020 15988
rect 573076 15932 573086 15988
rect 361172 15764 361228 15932
rect 361172 15708 367948 15764
rect 368004 15708 368014 15764
rect 117618 15036 117628 15092
rect 117684 15036 121884 15092
rect 121940 15036 121950 15092
rect 122770 15036 122780 15092
rect 122836 15036 126924 15092
rect 126980 15036 126990 15092
rect 120978 14924 120988 14980
rect 121044 14924 125020 14980
rect 125076 14924 125086 14980
rect 235442 14924 235452 14980
rect 235508 14924 253708 14980
rect 253764 14924 253774 14980
rect 126018 14812 126028 14868
rect 126084 14812 129724 14868
rect 129780 14812 129790 14868
rect 233874 14812 233884 14868
rect 233940 14812 252028 14868
rect 252084 14812 252094 14868
rect 119298 14700 119308 14756
rect 119364 14700 123452 14756
rect 123508 14700 123518 14756
rect 232306 14700 232316 14756
rect 232372 14700 250460 14756
rect 250516 14700 250526 14756
rect 422034 14700 422044 14756
rect 422100 14700 480508 14756
rect 480564 14700 480574 14756
rect 229170 14588 229180 14644
rect 229236 14588 246988 14644
rect 247044 14588 247054 14644
rect 359314 14588 359324 14644
rect 359380 14588 404908 14644
rect 404964 14588 404974 14644
rect 459666 14588 459676 14644
rect 459732 14588 525868 14644
rect 525924 14588 525934 14644
rect 227602 14476 227612 14532
rect 227668 14476 245532 14532
rect 245588 14476 245598 14532
rect 374098 14476 374108 14532
rect 374164 14476 389788 14532
rect 389844 14476 389854 14532
rect 390674 14476 390684 14532
rect 390740 14476 443548 14532
rect 443604 14476 443614 14532
rect 451826 14476 451836 14532
rect 451892 14476 517468 14532
rect 517524 14476 517534 14532
rect 124338 14364 124348 14420
rect 124404 14364 128156 14420
rect 128212 14364 128222 14420
rect 230738 14364 230748 14420
rect 230804 14364 248780 14420
rect 248836 14364 248846 14420
rect 275426 14364 275436 14420
rect 275492 14364 300748 14420
rect 300804 14364 300814 14420
rect 316642 14364 316652 14420
rect 316708 14364 349468 14420
rect 349524 14364 349534 14420
rect 352706 14364 352716 14420
rect 352772 14364 386540 14420
rect 386596 14364 386606 14420
rect 387986 14364 387996 14420
rect 388052 14364 396508 14420
rect 396564 14364 396574 14420
rect 404786 14364 404796 14420
rect 404852 14364 460348 14420
rect 460404 14364 460414 14420
rect 478482 14364 478492 14420
rect 478548 14364 549388 14420
rect 549444 14364 549454 14420
rect 31938 14252 31948 14308
rect 32004 14252 51324 14308
rect 51380 14252 51390 14308
rect 226034 14252 226044 14308
rect 226100 14252 243740 14308
rect 243796 14252 243806 14308
rect 296594 14252 296604 14308
rect 296660 14252 329308 14308
rect 329364 14252 329374 14308
rect 335346 14252 335356 14308
rect 335412 14252 373100 14308
rect 373156 14252 373166 14308
rect 378130 14252 378140 14308
rect 378196 14252 428428 14308
rect 428484 14252 428494 14308
rect 429874 14252 429884 14308
rect 429940 14252 490700 14308
rect 490756 14252 490766 14308
rect 504018 14252 504028 14308
rect 504084 14252 581308 14308
rect 581364 14252 581374 14308
rect 131282 13356 131292 13412
rect 131348 13356 132860 13412
rect 132916 13356 132926 13412
rect 134530 13356 134540 13412
rect 134596 13356 136108 13412
rect 136164 13356 136174 13412
rect 139458 13356 139468 13412
rect 139524 13356 141148 13412
rect 141204 13356 141214 13412
rect 72370 13244 72380 13300
rect 72436 13244 84252 13300
rect 84308 13244 84318 13300
rect 129378 13244 129388 13300
rect 129444 13244 131404 13300
rect 131460 13244 131470 13300
rect 132738 13244 132748 13300
rect 132804 13244 134428 13300
rect 134484 13244 134494 13300
rect 137890 13244 137900 13300
rect 137956 13244 139580 13300
rect 139636 13244 139646 13300
rect 74162 13132 74172 13188
rect 74228 13132 85820 13188
rect 85876 13132 85886 13188
rect 80658 13020 80668 13076
rect 80724 13020 92428 13076
rect 92484 13020 92494 13076
rect 383506 13020 383516 13076
rect 383572 13020 430220 13076
rect 430276 13020 430286 13076
rect 450370 13020 450380 13076
rect 450436 13020 502572 13076
rect 502628 13020 502638 13076
rect 82338 12908 82348 12964
rect 82404 12908 94220 12964
rect 94276 12908 94286 12964
rect 388882 12908 388892 12964
rect 388948 12908 425180 12964
rect 425236 12908 425246 12964
rect 427298 12908 427308 12964
rect 427364 12908 478828 12964
rect 478884 12908 478894 12964
rect 77298 12796 77308 12852
rect 77364 12796 89180 12852
rect 89236 12796 89246 12852
rect 346098 12796 346108 12852
rect 346164 12796 388108 12852
rect 388164 12796 388174 12852
rect 396946 12796 396956 12852
rect 397012 12796 450268 12852
rect 450324 12796 450334 12852
rect 469074 12796 469084 12852
rect 469140 12796 537628 12852
rect 537684 12796 537694 12852
rect 75618 12684 75628 12740
rect 75684 12684 87388 12740
rect 87444 12684 87454 12740
rect 277778 12684 277788 12740
rect 277844 12684 305788 12740
rect 305844 12684 305854 12740
rect 306898 12684 306908 12740
rect 306964 12684 322588 12740
rect 322644 12684 322654 12740
rect 337362 12684 337372 12740
rect 337428 12684 378028 12740
rect 378084 12684 378094 12740
rect 409490 12684 409500 12740
rect 409556 12684 465388 12740
rect 465444 12684 465454 12740
rect 483186 12684 483196 12740
rect 483252 12684 554428 12740
rect 554484 12684 554494 12740
rect 15138 12572 15148 12628
rect 15204 12572 37212 12628
rect 37268 12572 37278 12628
rect 78978 12572 78988 12628
rect 79044 12572 90972 12628
rect 91028 12572 91038 12628
rect 301298 12572 301308 12628
rect 301364 12572 334348 12628
rect 334404 12572 334414 12628
rect 362450 12572 362460 12628
rect 362516 12572 408268 12628
rect 408324 12572 408334 12628
rect 423602 12572 423612 12628
rect 423668 12572 482188 12628
rect 482244 12572 482254 12628
rect 484754 12572 484764 12628
rect 484820 12572 557788 12628
rect 557844 12572 557854 12628
rect 136098 12012 136108 12068
rect 136164 12012 138012 12068
rect 138068 12012 138078 12068
rect 45826 11564 45836 11620
rect 45892 11564 62300 11620
rect 62356 11564 62366 11620
rect 207218 11564 207228 11620
rect 207284 11564 220780 11620
rect 220836 11564 220846 11620
rect 49634 11452 49644 11508
rect 49700 11452 65660 11508
rect 65716 11452 65726 11508
rect 211922 11452 211932 11508
rect 211988 11452 226492 11508
rect 226548 11452 226558 11508
rect 55346 11340 55356 11396
rect 55412 11340 70588 11396
rect 70644 11340 70654 11396
rect 210354 11340 210364 11396
rect 210420 11340 224588 11396
rect 224644 11340 224654 11396
rect 412626 11340 412636 11396
rect 412692 11340 470204 11396
rect 470260 11340 470270 11396
rect 47730 11228 47740 11284
rect 47796 11228 63980 11284
rect 64036 11228 64046 11284
rect 204082 11228 204092 11284
rect 204148 11228 216972 11284
rect 217028 11228 217038 11284
rect 418898 11228 418908 11284
rect 418964 11228 477820 11284
rect 477876 11228 477886 11284
rect 51538 11116 51548 11172
rect 51604 11116 67452 11172
rect 67508 11116 67518 11172
rect 208786 11116 208796 11172
rect 208852 11116 222684 11172
rect 222740 11116 222750 11172
rect 349906 11116 349916 11172
rect 349972 11116 394044 11172
rect 394100 11116 394110 11172
rect 465938 11116 465948 11172
rect 466004 11116 534940 11172
rect 534996 11116 535006 11172
rect 43922 11004 43932 11060
rect 43988 11004 60732 11060
rect 60788 11004 60798 11060
rect 205650 11004 205660 11060
rect 205716 11004 218876 11060
rect 218932 11004 218942 11060
rect 312386 11004 312396 11060
rect 312452 11004 346444 11060
rect 346500 11004 346510 11060
rect 360882 11004 360892 11060
rect 360948 11004 407372 11060
rect 407428 11004 407438 11060
rect 407586 11004 407596 11060
rect 407652 11004 437836 11060
rect 437892 11004 437902 11060
rect 461234 11004 461244 11060
rect 461300 11004 529228 11060
rect 529284 11004 529294 11060
rect 531458 11004 531468 11060
rect 531524 11004 571228 11060
rect 571284 11004 571294 11060
rect 13346 10892 13356 10948
rect 13412 10892 35644 10948
rect 35700 10892 35710 10948
rect 53442 10892 53452 10948
rect 53508 10892 68908 10948
rect 68964 10892 68974 10948
rect 202514 10892 202524 10948
rect 202580 10892 215068 10948
rect 215124 10892 215134 10948
rect 299730 10892 299740 10948
rect 299796 10892 333116 10948
rect 333172 10892 333182 10948
rect 334226 10892 334236 10948
rect 334292 10892 361228 10948
rect 375666 10892 375676 10948
rect 375732 10892 424508 10948
rect 424564 10892 424574 10948
rect 433010 10892 433020 10948
rect 433076 10892 494956 10948
rect 495012 10892 495022 10948
rect 502292 10892 569212 10948
rect 569268 10892 569278 10948
rect 361172 10836 361228 10892
rect 502292 10836 502348 10892
rect 361172 10780 375004 10836
rect 375060 10780 375070 10836
rect 494162 10780 494172 10836
rect 494228 10780 502348 10836
rect 412066 9548 412076 9604
rect 412132 9548 464492 9604
rect 464548 9548 464558 9604
rect 365586 9436 365596 9492
rect 365652 9436 413084 9492
rect 413140 9436 413150 9492
rect 459218 9436 459228 9492
rect 459284 9436 514108 9492
rect 514164 9436 514174 9492
rect 320114 9324 320124 9380
rect 320180 9324 357868 9380
rect 357924 9324 357934 9380
rect 395378 9324 395388 9380
rect 395444 9324 449260 9380
rect 449316 9324 449326 9380
rect 480834 9324 480844 9380
rect 480900 9324 544460 9380
rect 544516 9324 544526 9380
rect 252690 9212 252700 9268
rect 252756 9212 275996 9268
rect 276052 9212 276062 9268
rect 306002 9212 306012 9268
rect 306068 9212 340732 9268
rect 340788 9212 340798 9268
rect 357746 9212 357756 9268
rect 357812 9212 403564 9268
rect 403620 9212 403630 9268
rect 406354 9212 406364 9268
rect 406420 9212 462588 9268
rect 462644 9212 462654 9268
rect 480050 9212 480060 9268
rect 480116 9212 552076 9268
rect 552132 9212 552142 9268
rect -960 8596 480 8792
rect -960 8568 8428 8596
rect 392 8540 8428 8568
rect 8372 8484 8428 8540
rect 8372 8428 530908 8484
rect 530964 8428 530974 8484
rect 360322 7980 360332 8036
rect 360388 7980 395948 8036
rect 396004 7980 396014 8036
rect 431732 7980 441644 8036
rect 441700 7980 441710 8036
rect 444322 7980 444332 8036
rect 444388 7980 458780 8036
rect 458836 7980 458846 8036
rect 478772 7980 498764 8036
rect 498820 7980 498830 8036
rect 431732 7924 431788 7980
rect 478772 7924 478828 7980
rect 289762 7868 289772 7924
rect 289828 7868 304556 7924
rect 304612 7868 304622 7924
rect 337698 7868 337708 7924
rect 337764 7868 380716 7924
rect 380772 7868 380782 7924
rect 388210 7868 388220 7924
rect 388276 7868 431788 7924
rect 440962 7868 440972 7924
rect 441028 7868 478828 7924
rect 491372 7868 496860 7924
rect 496916 7868 496926 7924
rect 498082 7868 498092 7924
rect 498148 7868 525420 7924
rect 525476 7868 525486 7924
rect 491372 7812 491428 7868
rect 261202 7756 261212 7812
rect 261268 7756 281708 7812
rect 281764 7756 281774 7812
rect 296482 7756 296492 7812
rect 296548 7756 327404 7812
rect 327460 7756 327470 7812
rect 341058 7756 341068 7812
rect 341124 7756 384524 7812
rect 384580 7756 384590 7812
rect 433458 7756 433468 7812
rect 433524 7756 491428 7812
rect 496402 7756 496412 7812
rect 496468 7756 553980 7812
rect 554036 7756 554046 7812
rect 265458 7644 265468 7700
rect 265524 7644 293132 7700
rect 293188 7644 293198 7700
rect 304098 7644 304108 7700
rect 304164 7644 338828 7700
rect 338884 7644 338894 7700
rect 379698 7644 379708 7700
rect 379764 7644 432124 7700
rect 432180 7644 432190 7700
rect 445330 7644 445340 7700
rect 445396 7644 510188 7700
rect 510244 7644 510254 7700
rect 548482 7644 548492 7700
rect 548548 7644 580636 7700
rect 580692 7644 580702 7700
rect 11554 7532 11564 7588
rect 11620 7532 33740 7588
rect 33796 7532 33806 7588
rect 247090 7532 247100 7588
rect 247156 7532 270284 7588
rect 270340 7532 270350 7588
rect 280578 7532 280588 7588
rect 280644 7532 307580 7588
rect 307636 7532 307646 7588
rect 322690 7532 322700 7588
rect 322756 7532 361676 7588
rect 361732 7532 361742 7588
rect 383058 7532 383068 7588
rect 383124 7532 435932 7588
rect 435988 7532 435998 7588
rect 436818 7532 436828 7588
rect 436884 7532 500668 7588
rect 500724 7532 500734 7588
rect 506482 7532 506492 7588
rect 506548 7532 567308 7588
rect 567364 7532 567374 7588
rect 594514 7308 594524 7364
rect 594580 7336 595672 7364
rect 594580 7308 597000 7336
rect 595560 7112 597000 7308
rect 314962 6748 314972 6804
rect 315028 6748 321692 6804
rect 321748 6748 321758 6804
rect 456082 6636 456092 6692
rect 456148 6636 456988 6692
rect 457044 6636 457054 6692
rect 176418 6412 176428 6468
rect 176484 6412 184604 6468
rect 184660 6412 184670 6468
rect 191650 6412 191660 6468
rect 191716 6412 203644 6468
rect 203700 6412 203710 6468
rect 400642 6412 400652 6468
rect 400708 6412 434028 6468
rect 434084 6412 434094 6468
rect 186498 6300 186508 6356
rect 186564 6300 196028 6356
rect 196084 6300 196094 6356
rect 196578 6300 196588 6356
rect 196644 6300 209356 6356
rect 209412 6300 209422 6356
rect 346882 6300 346892 6356
rect 346948 6300 365484 6356
rect 365540 6300 365550 6356
rect 393138 6300 393148 6356
rect 393204 6300 447356 6356
rect 447412 6300 447422 6356
rect 467842 6300 467852 6356
rect 467908 6300 508284 6356
rect 508340 6300 508350 6356
rect 174738 6188 174748 6244
rect 174804 6188 182700 6244
rect 182756 6188 182766 6244
rect 183138 6188 183148 6244
rect 183204 6188 192220 6244
rect 192276 6188 192286 6244
rect 194898 6188 194908 6244
rect 194964 6188 207452 6244
rect 207508 6188 207518 6244
rect 308242 6188 308252 6244
rect 308308 6188 319788 6244
rect 319844 6188 319854 6244
rect 336802 6188 336812 6244
rect 336868 6188 344540 6244
rect 344596 6188 344606 6244
rect 353602 6188 353612 6244
rect 353668 6188 376908 6244
rect 376964 6188 376974 6244
rect 419122 6188 419132 6244
rect 419188 6188 474012 6244
rect 474068 6188 474078 6244
rect 477922 6188 477932 6244
rect 477988 6188 487340 6244
rect 487396 6188 487406 6244
rect 501442 6188 501452 6244
rect 501508 6188 515900 6244
rect 515956 6188 515966 6244
rect 171378 6076 171388 6132
rect 171444 6076 178892 6132
rect 178948 6076 178958 6132
rect 181458 6076 181468 6132
rect 181524 6076 190316 6132
rect 190372 6076 190382 6132
rect 198258 6076 198268 6132
rect 198324 6076 211260 6132
rect 211316 6076 211326 6132
rect 241938 6076 241948 6132
rect 242004 6076 264572 6132
rect 264628 6076 264638 6132
rect 317538 6076 317548 6132
rect 317604 6076 355964 6132
rect 356020 6076 356030 6132
rect 377122 6076 377132 6132
rect 377188 6076 401660 6132
rect 401716 6076 401726 6132
rect 430098 6076 430108 6132
rect 430164 6076 493052 6132
rect 493108 6076 493118 6132
rect 503122 6076 503132 6132
rect 503188 6076 533036 6132
rect 533092 6076 533102 6132
rect 168130 5964 168140 6020
rect 168196 5964 175084 6020
rect 175140 5964 175150 6020
rect 188178 5964 188188 6020
rect 188244 5964 188692 6020
rect 193218 5964 193228 6020
rect 193284 5964 205548 6020
rect 205604 5964 205614 6020
rect 215170 5964 215180 6020
rect 215236 5964 230300 6020
rect 230356 5964 230366 6020
rect 253810 5964 253820 6020
rect 253876 5964 277900 6020
rect 277956 5964 277966 6020
rect 283938 5964 283948 6020
rect 284004 5964 314188 6020
rect 314244 5964 314254 6020
rect 327618 5964 327628 6020
rect 327684 5964 367388 6020
rect 367444 5964 367454 6020
rect 369618 5964 369628 6020
rect 369684 5964 418796 6020
rect 418852 5964 418862 6020
rect 456194 5964 456204 6020
rect 456260 5964 512092 6020
rect 512148 5964 512158 6020
rect 513202 5964 513212 6020
rect 513268 5964 574924 6020
rect 574980 5964 574990 6020
rect 188636 5908 188692 5964
rect 22978 5852 22988 5908
rect 23044 5852 32732 5908
rect 32788 5852 32798 5908
rect 169698 5852 169708 5908
rect 169764 5852 176988 5908
rect 177044 5852 177054 5908
rect 179778 5852 179788 5908
rect 179844 5852 188412 5908
rect 188468 5852 188478 5908
rect 188636 5852 197932 5908
rect 197988 5852 197998 5908
rect 199938 5852 199948 5908
rect 200004 5852 213164 5908
rect 213220 5852 213230 5908
rect 213378 5852 213388 5908
rect 213444 5852 228508 5908
rect 228564 5852 228574 5908
rect 262098 5852 262108 5908
rect 262164 5852 289324 5908
rect 289380 5852 289390 5908
rect 292338 5852 292348 5908
rect 292404 5852 325500 5908
rect 325556 5852 325566 5908
rect 343522 5852 343532 5908
rect 343588 5852 354060 5908
rect 354116 5852 354126 5908
rect 354498 5852 354508 5908
rect 354564 5852 399868 5908
rect 399924 5852 399934 5908
rect 413298 5852 413308 5908
rect 413364 5852 448812 5908
rect 448868 5852 448878 5908
rect 456306 5852 456316 5908
rect 456372 5852 472108 5908
rect 472164 5852 472174 5908
rect 487218 5852 487228 5908
rect 487284 5852 561036 5908
rect 561092 5852 561102 5908
rect 178098 5740 178108 5796
rect 178164 5740 186508 5796
rect 186564 5740 186574 5796
rect 414082 5404 414092 5460
rect 414148 5404 416892 5460
rect 416948 5404 416958 5460
rect 173058 5068 173068 5124
rect 173124 5068 180796 5124
rect 180852 5068 180862 5124
rect 184818 5068 184828 5124
rect 184884 5068 194124 5124
rect 194180 5068 194190 5124
rect 449362 5068 449372 5124
rect 449428 5068 453068 5124
rect 453124 5068 453134 5124
rect 147858 4956 147868 5012
rect 147924 4956 150332 5012
rect 150388 4956 150398 5012
rect 278898 4956 278908 5012
rect 278964 4956 308364 5012
rect 308420 4956 308430 5012
rect 159618 4844 159628 4900
rect 159684 4844 163660 4900
rect 163716 4844 163726 4900
rect 282258 4844 282268 4900
rect 282324 4844 312172 4900
rect 312228 4844 312238 4900
rect 467058 4844 467068 4900
rect 467124 4844 536844 4900
rect 536900 4844 536910 4900
rect 158050 4732 158060 4788
rect 158116 4732 161756 4788
rect 161812 4732 161822 4788
rect 168018 4732 168028 4788
rect 168084 4732 173180 4788
rect 173236 4732 173246 4788
rect 250338 4732 250348 4788
rect 250404 4732 274092 4788
rect 274148 4732 274158 4788
rect 297490 4732 297500 4788
rect 297556 4732 331212 4788
rect 331268 4732 331278 4788
rect 462018 4732 462028 4788
rect 462084 4732 531132 4788
rect 531188 4732 531198 4788
rect 577042 4732 577052 4788
rect 577108 4732 584444 4788
rect 584500 4732 584510 4788
rect 28690 4620 28700 4676
rect 28756 4620 48748 4676
rect 48804 4620 48814 4676
rect 144722 4620 144732 4676
rect 144788 4620 146524 4676
rect 146580 4620 146590 4676
rect 154578 4620 154588 4676
rect 154644 4620 157948 4676
rect 158004 4620 158014 4676
rect 237010 4620 237020 4676
rect 237076 4620 257068 4676
rect 257124 4620 257134 4676
rect 267250 4620 267260 4676
rect 267316 4620 295036 4676
rect 295092 4620 295102 4676
rect 307458 4620 307468 4676
rect 307524 4620 342748 4676
rect 342804 4620 342814 4676
rect 472210 4620 472220 4676
rect 472276 4620 542668 4676
rect 542724 4620 542734 4676
rect 24882 4508 24892 4564
rect 24948 4508 45388 4564
rect 45444 4508 45454 4564
rect 166338 4508 166348 4564
rect 166404 4508 171388 4564
rect 171444 4508 171454 4564
rect 240370 4508 240380 4564
rect 240436 4508 262668 4564
rect 262724 4508 262734 4564
rect 263778 4508 263788 4564
rect 263844 4508 291228 4564
rect 291284 4508 291294 4564
rect 307570 4508 307580 4564
rect 307636 4508 310268 4564
rect 310324 4508 310334 4564
rect 310818 4508 310828 4564
rect 310884 4508 348348 4564
rect 348404 4508 348414 4564
rect 475570 4508 475580 4564
rect 475636 4508 548268 4564
rect 548324 4508 548334 4564
rect 26786 4396 26796 4452
rect 26852 4396 47068 4452
rect 47124 4396 47134 4452
rect 238690 4396 238700 4452
rect 238756 4396 260764 4452
rect 260820 4396 260830 4452
rect 273858 4396 273868 4452
rect 273924 4396 302652 4452
rect 302708 4396 302718 4452
rect 320898 4396 320908 4452
rect 320964 4396 359772 4452
rect 359828 4396 359838 4452
rect 485538 4396 485548 4452
rect 485604 4396 559692 4452
rect 559748 4396 559758 4452
rect 21074 4284 21084 4340
rect 21140 4284 42028 4340
rect 42084 4284 42094 4340
rect 57250 4284 57260 4340
rect 57316 4284 72268 4340
rect 72324 4284 72334 4340
rect 146178 4284 146188 4340
rect 146244 4284 148428 4340
rect 148484 4284 148494 4340
rect 149538 4284 149548 4340
rect 149604 4284 152236 4340
rect 152292 4284 152302 4340
rect 152898 4284 152908 4340
rect 152964 4284 156044 4340
rect 156100 4284 156110 4340
rect 162978 4284 162988 4340
rect 163044 4284 167468 4340
rect 167524 4284 167534 4340
rect 191538 4284 191548 4340
rect 191604 4284 201740 4340
rect 201796 4284 201806 4340
rect 248658 4284 248668 4340
rect 248724 4284 272188 4340
rect 272244 4284 272254 4340
rect 285730 4284 285740 4340
rect 285796 4284 317884 4340
rect 317940 4284 317950 4340
rect 330978 4284 330988 4340
rect 331044 4284 371308 4340
rect 371364 4284 371374 4340
rect 490578 4284 490588 4340
rect 490644 4284 565404 4340
rect 565460 4284 565470 4340
rect 17266 4172 17276 4228
rect 17332 4172 38780 4228
rect 38836 4172 38846 4228
rect 59154 4172 59164 4228
rect 59220 4172 74284 4228
rect 74340 4172 74350 4228
rect 151218 4172 151228 4228
rect 151284 4172 154140 4228
rect 154196 4172 154206 4228
rect 156258 4172 156268 4228
rect 156324 4172 159852 4228
rect 159908 4172 159918 4228
rect 161298 4172 161308 4228
rect 161364 4172 165564 4228
rect 165620 4172 165630 4228
rect 189858 4172 189868 4228
rect 189924 4172 199948 4228
rect 200004 4172 200014 4228
rect 257842 4172 257852 4228
rect 257908 4172 258860 4228
rect 258916 4172 258926 4228
rect 268818 4172 268828 4228
rect 268884 4172 296940 4228
rect 296996 4172 297006 4228
rect 302418 4172 302428 4228
rect 302484 4172 336924 4228
rect 336980 4172 336990 4228
rect 339378 4172 339388 4228
rect 339444 4172 382620 4228
rect 382676 4172 382686 4228
rect 498978 4172 498988 4228
rect 499044 4172 576828 4228
rect 576884 4172 576894 4228
rect 164658 4060 164668 4116
rect 164724 4060 169372 4116
rect 169428 4060 169438 4116
rect 243618 4060 243628 4116
rect 243684 4060 266476 4116
rect 266532 4060 266542 4116
rect 266700 4060 283612 4116
rect 283668 4060 283678 4116
rect 266700 4004 266756 4060
rect 258738 3948 258748 4004
rect 258804 3948 266756 4004
rect 267092 3948 279804 4004
rect 279860 3948 279870 4004
rect 267092 3892 267148 3948
rect 255378 3836 255388 3892
rect 255444 3836 267148 3892
rect 365362 2940 365372 2996
rect 365428 2940 411180 2996
rect 411236 2940 411246 2996
rect 464594 2828 464604 2884
rect 464660 2828 519708 2884
rect 519764 2828 519774 2884
rect 409938 2716 409948 2772
rect 410004 2716 468300 2772
rect 468356 2716 468366 2772
rect 484642 2716 484652 2772
rect 484708 2716 546364 2772
rect 546420 2716 546430 2772
rect 371410 2604 371420 2660
rect 371476 2604 420700 2660
rect 420756 2604 420766 2660
rect 426738 2604 426748 2660
rect 426804 2604 489244 2660
rect 489300 2604 489310 2660
rect 324258 2492 324268 2548
rect 324324 2492 363580 2548
rect 363636 2492 363646 2548
rect 386418 2492 386428 2548
rect 386484 2492 439740 2548
rect 439796 2492 439806 2548
rect 441858 2492 441868 2548
rect 441924 2492 506380 2548
rect 506436 2492 506446 2548
rect 425394 28 425404 84
rect 425460 28 485772 84
rect 485828 28 485838 84
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 3154 597212 3774 598268
rect 3154 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 3774 597212
rect 3154 597088 3774 597156
rect 3154 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 3774 597088
rect 3154 596964 3774 597032
rect 3154 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 3774 596964
rect 3154 596840 3774 596908
rect 3154 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 3774 596840
rect 3154 580350 3774 596784
rect 3154 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 3774 580350
rect 3154 580226 3774 580294
rect 3154 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 3774 580226
rect 3154 580102 3774 580170
rect 3154 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 3774 580102
rect 3154 579978 3774 580046
rect 3154 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 3774 579978
rect 3154 562350 3774 579922
rect 3154 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 3774 562350
rect 3154 562226 3774 562294
rect 3154 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 3774 562226
rect 3154 562102 3774 562170
rect 3154 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 3774 562102
rect 3154 561978 3774 562046
rect 3154 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 3774 561978
rect 3154 544350 3774 561922
rect 3154 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 3774 544350
rect 3154 544226 3774 544294
rect 3154 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 3774 544226
rect 3154 544102 3774 544170
rect 3154 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 3774 544102
rect 3154 543978 3774 544046
rect 3154 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 3774 543978
rect 3154 526350 3774 543922
rect 3154 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 3774 526350
rect 3154 526226 3774 526294
rect 3154 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 3774 526226
rect 3154 526102 3774 526170
rect 3154 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 3774 526102
rect 3154 525978 3774 526046
rect 3154 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 3774 525978
rect 3154 508350 3774 525922
rect 3154 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 3774 508350
rect 3154 508226 3774 508294
rect 3154 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 3774 508226
rect 3154 508102 3774 508170
rect 3154 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 3774 508102
rect 3154 507978 3774 508046
rect 3154 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 3774 507978
rect 3154 490350 3774 507922
rect 3154 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 3774 490350
rect 3154 490226 3774 490294
rect 3154 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 3774 490226
rect 3154 490102 3774 490170
rect 3154 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 3774 490102
rect 3154 489978 3774 490046
rect 3154 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 3774 489978
rect 3154 472350 3774 489922
rect 3154 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 3774 472350
rect 3154 472226 3774 472294
rect 3154 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 3774 472226
rect 3154 472102 3774 472170
rect 3154 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 3774 472102
rect 3154 471978 3774 472046
rect 3154 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 3774 471978
rect 3154 454350 3774 471922
rect 3154 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 3774 454350
rect 3154 454226 3774 454294
rect 3154 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 3774 454226
rect 3154 454102 3774 454170
rect 3154 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 3774 454102
rect 3154 453978 3774 454046
rect 3154 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 3774 453978
rect 3154 436350 3774 453922
rect 3154 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 3774 436350
rect 3154 436226 3774 436294
rect 3154 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 3774 436226
rect 3154 436102 3774 436170
rect 3154 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 3774 436102
rect 3154 435978 3774 436046
rect 3154 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 3774 435978
rect 3154 418350 3774 435922
rect 3154 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 3774 418350
rect 3154 418226 3774 418294
rect 3154 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 3774 418226
rect 3154 418102 3774 418170
rect 3154 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 3774 418102
rect 3154 417978 3774 418046
rect 3154 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 3774 417978
rect 3154 400350 3774 417922
rect 3154 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 3774 400350
rect 3154 400226 3774 400294
rect 3154 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 3774 400226
rect 3154 400102 3774 400170
rect 3154 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 3774 400102
rect 3154 399978 3774 400046
rect 3154 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 3774 399978
rect 3154 382350 3774 399922
rect 3154 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 3774 382350
rect 3154 382226 3774 382294
rect 3154 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 3774 382226
rect 3154 382102 3774 382170
rect 3154 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 3774 382102
rect 3154 381978 3774 382046
rect 3154 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 3774 381978
rect 3154 364350 3774 381922
rect 3154 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 3774 364350
rect 3154 364226 3774 364294
rect 3154 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 3774 364226
rect 3154 364102 3774 364170
rect 3154 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 3774 364102
rect 3154 363978 3774 364046
rect 3154 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 3774 363978
rect 3154 346350 3774 363922
rect 3154 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 3774 346350
rect 3154 346226 3774 346294
rect 3154 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 3774 346226
rect 3154 346102 3774 346170
rect 3154 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 3774 346102
rect 3154 345978 3774 346046
rect 3154 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 3774 345978
rect 3154 328350 3774 345922
rect 3154 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 3774 328350
rect 3154 328226 3774 328294
rect 3154 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 3774 328226
rect 3154 328102 3774 328170
rect 3154 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 3774 328102
rect 3154 327978 3774 328046
rect 3154 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 3774 327978
rect 3154 310350 3774 327922
rect 3154 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 3774 310350
rect 3154 310226 3774 310294
rect 3154 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 3774 310226
rect 3154 310102 3774 310170
rect 3154 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 3774 310102
rect 3154 309978 3774 310046
rect 3154 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 3774 309978
rect 3154 292350 3774 309922
rect 3154 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 3774 292350
rect 3154 292226 3774 292294
rect 3154 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 3774 292226
rect 3154 292102 3774 292170
rect 3154 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 3774 292102
rect 3154 291978 3774 292046
rect 3154 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 3774 291978
rect 3154 274350 3774 291922
rect 3154 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 3774 274350
rect 3154 274226 3774 274294
rect 3154 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 3774 274226
rect 3154 274102 3774 274170
rect 3154 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 3774 274102
rect 3154 273978 3774 274046
rect 3154 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 3774 273978
rect 3154 256350 3774 273922
rect 3154 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 3774 256350
rect 3154 256226 3774 256294
rect 3154 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 3774 256226
rect 3154 256102 3774 256170
rect 3154 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 3774 256102
rect 3154 255978 3774 256046
rect 3154 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 3774 255978
rect 3154 238350 3774 255922
rect 3154 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 3774 238350
rect 3154 238226 3774 238294
rect 3154 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 3774 238226
rect 3154 238102 3774 238170
rect 3154 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 3774 238102
rect 3154 237978 3774 238046
rect 3154 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 3774 237978
rect 3154 220350 3774 237922
rect 3154 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 3774 220350
rect 3154 220226 3774 220294
rect 3154 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 3774 220226
rect 3154 220102 3774 220170
rect 3154 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 3774 220102
rect 3154 219978 3774 220046
rect 3154 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 3774 219978
rect 3154 202350 3774 219922
rect 3154 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 3774 202350
rect 3154 202226 3774 202294
rect 3154 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 3774 202226
rect 3154 202102 3774 202170
rect 3154 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 3774 202102
rect 3154 201978 3774 202046
rect 3154 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 3774 201978
rect 3154 184350 3774 201922
rect 3154 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 3774 184350
rect 3154 184226 3774 184294
rect 3154 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 3774 184226
rect 3154 184102 3774 184170
rect 3154 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 3774 184102
rect 3154 183978 3774 184046
rect 3154 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 3774 183978
rect 3154 166350 3774 183922
rect 3154 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 3774 166350
rect 3154 166226 3774 166294
rect 3154 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 3774 166226
rect 3154 166102 3774 166170
rect 3154 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 3774 166102
rect 3154 165978 3774 166046
rect 3154 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 3774 165978
rect 3154 148350 3774 165922
rect 3154 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 3774 148350
rect 3154 148226 3774 148294
rect 3154 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 3774 148226
rect 3154 148102 3774 148170
rect 3154 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 3774 148102
rect 3154 147978 3774 148046
rect 3154 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 3774 147978
rect 3154 130350 3774 147922
rect 3154 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 3774 130350
rect 3154 130226 3774 130294
rect 3154 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 3774 130226
rect 3154 130102 3774 130170
rect 3154 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 3774 130102
rect 3154 129978 3774 130046
rect 3154 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 3774 129978
rect 3154 112350 3774 129922
rect 3154 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 3774 112350
rect 3154 112226 3774 112294
rect 3154 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 3774 112226
rect 3154 112102 3774 112170
rect 3154 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 3774 112102
rect 3154 111978 3774 112046
rect 3154 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 3774 111978
rect 3154 94350 3774 111922
rect 3154 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 3774 94350
rect 3154 94226 3774 94294
rect 3154 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 3774 94226
rect 3154 94102 3774 94170
rect 3154 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 3774 94102
rect 3154 93978 3774 94046
rect 3154 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 3774 93978
rect 3154 76350 3774 93922
rect 3154 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 3774 76350
rect 3154 76226 3774 76294
rect 3154 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 3774 76226
rect 3154 76102 3774 76170
rect 3154 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 3774 76102
rect 3154 75978 3774 76046
rect 3154 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 3774 75978
rect 3154 58350 3774 75922
rect 3154 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 3774 58350
rect 3154 58226 3774 58294
rect 3154 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 3774 58226
rect 3154 58102 3774 58170
rect 3154 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 3774 58102
rect 3154 57978 3774 58046
rect 3154 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 3774 57978
rect 3154 40350 3774 57922
rect 3154 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 3774 40350
rect 3154 40226 3774 40294
rect 3154 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 3774 40226
rect 3154 40102 3774 40170
rect 3154 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 3774 40102
rect 3154 39978 3774 40046
rect 3154 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 3774 39978
rect 3154 22350 3774 39922
rect 3154 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 3774 22350
rect 3154 22226 3774 22294
rect 3154 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 3774 22226
rect 3154 22102 3774 22170
rect 3154 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 3774 22102
rect 3154 21978 3774 22046
rect 3154 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 3774 21978
rect 3154 4350 3774 21922
rect 3154 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 3774 4350
rect 3154 4226 3774 4294
rect 3154 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 3774 4226
rect 3154 4102 3774 4170
rect 3154 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 3774 4102
rect 3154 3978 3774 4046
rect 3154 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 3774 3978
rect 3154 -160 3774 3922
rect 3154 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 3774 -160
rect 3154 -284 3774 -216
rect 3154 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 3774 -284
rect 3154 -408 3774 -340
rect 3154 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 3774 -408
rect 3154 -532 3774 -464
rect 3154 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 3774 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 3154 -1644 3774 -588
rect 6874 598172 7494 598268
rect 6874 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 7494 598172
rect 6874 598048 7494 598116
rect 6874 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 7494 598048
rect 6874 597924 7494 597992
rect 6874 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 7494 597924
rect 6874 597800 7494 597868
rect 6874 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 7494 597800
rect 6874 586350 7494 597744
rect 6874 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 7494 586350
rect 6874 586226 7494 586294
rect 6874 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 7494 586226
rect 6874 586102 7494 586170
rect 6874 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 7494 586102
rect 6874 585978 7494 586046
rect 6874 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 7494 585978
rect 6874 568350 7494 585922
rect 6874 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 7494 568350
rect 6874 568226 7494 568294
rect 6874 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 7494 568226
rect 6874 568102 7494 568170
rect 6874 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 7494 568102
rect 6874 567978 7494 568046
rect 6874 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 7494 567978
rect 6874 550350 7494 567922
rect 6874 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 7494 550350
rect 6874 550226 7494 550294
rect 6874 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 7494 550226
rect 6874 550102 7494 550170
rect 6874 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 7494 550102
rect 6874 549978 7494 550046
rect 6874 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 7494 549978
rect 6874 532350 7494 549922
rect 6874 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 7494 532350
rect 6874 532226 7494 532294
rect 6874 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 7494 532226
rect 6874 532102 7494 532170
rect 6874 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 7494 532102
rect 6874 531978 7494 532046
rect 6874 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 7494 531978
rect 6874 514350 7494 531922
rect 21154 597212 21774 598268
rect 21154 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 21774 597212
rect 21154 597088 21774 597156
rect 21154 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 21774 597088
rect 21154 596964 21774 597032
rect 21154 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 21774 596964
rect 21154 596840 21774 596908
rect 21154 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 21774 596840
rect 21154 580350 21774 596784
rect 21154 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 21774 580350
rect 21154 580226 21774 580294
rect 21154 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 21774 580226
rect 21154 580102 21774 580170
rect 21154 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 21774 580102
rect 21154 579978 21774 580046
rect 21154 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 21774 579978
rect 21154 562350 21774 579922
rect 21154 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 21774 562350
rect 21154 562226 21774 562294
rect 21154 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 21774 562226
rect 21154 562102 21774 562170
rect 21154 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 21774 562102
rect 21154 561978 21774 562046
rect 21154 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 21774 561978
rect 21154 544350 21774 561922
rect 21154 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 21774 544350
rect 21154 544226 21774 544294
rect 21154 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 21774 544226
rect 21154 544102 21774 544170
rect 21154 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 21774 544102
rect 21154 543978 21774 544046
rect 21154 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 21774 543978
rect 21154 526350 21774 543922
rect 21154 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 21774 526350
rect 21154 526226 21774 526294
rect 21154 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 21774 526226
rect 21154 526102 21774 526170
rect 21154 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 21774 526102
rect 21154 525978 21774 526046
rect 21154 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 21774 525978
rect 21154 520886 21774 525922
rect 24874 598172 25494 598268
rect 24874 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 25494 598172
rect 24874 598048 25494 598116
rect 24874 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 25494 598048
rect 24874 597924 25494 597992
rect 24874 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 25494 597924
rect 24874 597800 25494 597868
rect 24874 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 25494 597800
rect 24874 586350 25494 597744
rect 24874 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 25494 586350
rect 24874 586226 25494 586294
rect 24874 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 25494 586226
rect 24874 586102 25494 586170
rect 24874 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 25494 586102
rect 24874 585978 25494 586046
rect 24874 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 25494 585978
rect 24874 568350 25494 585922
rect 24874 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 25494 568350
rect 24874 568226 25494 568294
rect 24874 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 25494 568226
rect 24874 568102 25494 568170
rect 24874 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 25494 568102
rect 24874 567978 25494 568046
rect 24874 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 25494 567978
rect 24874 550350 25494 567922
rect 24874 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 25494 550350
rect 24874 550226 25494 550294
rect 24874 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 25494 550226
rect 24874 550102 25494 550170
rect 24874 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 25494 550102
rect 24874 549978 25494 550046
rect 24874 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 25494 549978
rect 24874 532350 25494 549922
rect 24874 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 25494 532350
rect 24874 532226 25494 532294
rect 24874 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 25494 532226
rect 24874 532102 25494 532170
rect 24874 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 25494 532102
rect 24874 531978 25494 532046
rect 24874 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 25494 531978
rect 24874 520886 25494 531922
rect 39154 597212 39774 598268
rect 39154 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 39774 597212
rect 39154 597088 39774 597156
rect 39154 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 39774 597088
rect 39154 596964 39774 597032
rect 39154 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 39774 596964
rect 39154 596840 39774 596908
rect 39154 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 39774 596840
rect 39154 580350 39774 596784
rect 39154 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 39774 580350
rect 39154 580226 39774 580294
rect 39154 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 39774 580226
rect 39154 580102 39774 580170
rect 39154 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 39774 580102
rect 39154 579978 39774 580046
rect 39154 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 39774 579978
rect 39154 562350 39774 579922
rect 39154 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 39774 562350
rect 39154 562226 39774 562294
rect 39154 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 39774 562226
rect 39154 562102 39774 562170
rect 39154 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 39774 562102
rect 39154 561978 39774 562046
rect 39154 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 39774 561978
rect 39154 544350 39774 561922
rect 39154 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 39774 544350
rect 39154 544226 39774 544294
rect 39154 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 39774 544226
rect 39154 544102 39774 544170
rect 39154 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 39774 544102
rect 39154 543978 39774 544046
rect 39154 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 39774 543978
rect 39154 526350 39774 543922
rect 39154 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 39774 526350
rect 39154 526226 39774 526294
rect 39154 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 39774 526226
rect 39154 526102 39774 526170
rect 39154 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 39774 526102
rect 39154 525978 39774 526046
rect 39154 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 39774 525978
rect 39154 520886 39774 525922
rect 42874 598172 43494 598268
rect 42874 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 43494 598172
rect 42874 598048 43494 598116
rect 42874 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 43494 598048
rect 42874 597924 43494 597992
rect 42874 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 43494 597924
rect 42874 597800 43494 597868
rect 42874 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 43494 597800
rect 42874 586350 43494 597744
rect 42874 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 43494 586350
rect 42874 586226 43494 586294
rect 42874 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 43494 586226
rect 42874 586102 43494 586170
rect 42874 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 43494 586102
rect 42874 585978 43494 586046
rect 42874 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 43494 585978
rect 42874 568350 43494 585922
rect 42874 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 43494 568350
rect 42874 568226 43494 568294
rect 42874 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 43494 568226
rect 42874 568102 43494 568170
rect 42874 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 43494 568102
rect 42874 567978 43494 568046
rect 42874 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 43494 567978
rect 42874 550350 43494 567922
rect 42874 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 43494 550350
rect 42874 550226 43494 550294
rect 42874 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 43494 550226
rect 42874 550102 43494 550170
rect 42874 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 43494 550102
rect 42874 549978 43494 550046
rect 42874 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 43494 549978
rect 42874 532350 43494 549922
rect 42874 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 43494 532350
rect 42874 532226 43494 532294
rect 42874 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 43494 532226
rect 42874 532102 43494 532170
rect 42874 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 43494 532102
rect 42874 531978 43494 532046
rect 42874 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 43494 531978
rect 42874 520886 43494 531922
rect 57154 597212 57774 598268
rect 57154 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 57774 597212
rect 57154 597088 57774 597156
rect 57154 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 57774 597088
rect 57154 596964 57774 597032
rect 57154 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 57774 596964
rect 57154 596840 57774 596908
rect 57154 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 57774 596840
rect 57154 580350 57774 596784
rect 57154 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 57774 580350
rect 57154 580226 57774 580294
rect 57154 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 57774 580226
rect 57154 580102 57774 580170
rect 57154 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 57774 580102
rect 57154 579978 57774 580046
rect 57154 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 57774 579978
rect 57154 562350 57774 579922
rect 57154 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 57774 562350
rect 57154 562226 57774 562294
rect 57154 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 57774 562226
rect 57154 562102 57774 562170
rect 57154 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 57774 562102
rect 57154 561978 57774 562046
rect 57154 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 57774 561978
rect 57154 544350 57774 561922
rect 57154 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 57774 544350
rect 57154 544226 57774 544294
rect 57154 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 57774 544226
rect 57154 544102 57774 544170
rect 57154 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 57774 544102
rect 57154 543978 57774 544046
rect 57154 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 57774 543978
rect 57154 526350 57774 543922
rect 57154 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 57774 526350
rect 57154 526226 57774 526294
rect 57154 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 57774 526226
rect 57154 526102 57774 526170
rect 57154 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 57774 526102
rect 57154 525978 57774 526046
rect 57154 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 57774 525978
rect 57154 520886 57774 525922
rect 60874 598172 61494 598268
rect 60874 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 61494 598172
rect 60874 598048 61494 598116
rect 60874 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 61494 598048
rect 60874 597924 61494 597992
rect 60874 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 61494 597924
rect 60874 597800 61494 597868
rect 60874 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 61494 597800
rect 60874 586350 61494 597744
rect 60874 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 61494 586350
rect 60874 586226 61494 586294
rect 60874 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 61494 586226
rect 60874 586102 61494 586170
rect 60874 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 61494 586102
rect 60874 585978 61494 586046
rect 60874 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 61494 585978
rect 60874 568350 61494 585922
rect 60874 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 61494 568350
rect 60874 568226 61494 568294
rect 60874 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 61494 568226
rect 60874 568102 61494 568170
rect 60874 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 61494 568102
rect 60874 567978 61494 568046
rect 60874 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 61494 567978
rect 60874 550350 61494 567922
rect 60874 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 61494 550350
rect 60874 550226 61494 550294
rect 60874 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 61494 550226
rect 60874 550102 61494 550170
rect 60874 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 61494 550102
rect 60874 549978 61494 550046
rect 60874 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 61494 549978
rect 60874 532350 61494 549922
rect 60874 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 61494 532350
rect 60874 532226 61494 532294
rect 60874 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 61494 532226
rect 60874 532102 61494 532170
rect 60874 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 61494 532102
rect 60874 531978 61494 532046
rect 60874 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 61494 531978
rect 60874 520886 61494 531922
rect 75154 597212 75774 598268
rect 75154 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 75774 597212
rect 75154 597088 75774 597156
rect 75154 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 75774 597088
rect 75154 596964 75774 597032
rect 75154 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 75774 596964
rect 75154 596840 75774 596908
rect 75154 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 75774 596840
rect 75154 580350 75774 596784
rect 75154 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 75774 580350
rect 75154 580226 75774 580294
rect 75154 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 75774 580226
rect 75154 580102 75774 580170
rect 75154 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 75774 580102
rect 75154 579978 75774 580046
rect 75154 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 75774 579978
rect 75154 562350 75774 579922
rect 75154 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 75774 562350
rect 75154 562226 75774 562294
rect 75154 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 75774 562226
rect 75154 562102 75774 562170
rect 75154 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 75774 562102
rect 75154 561978 75774 562046
rect 75154 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 75774 561978
rect 75154 544350 75774 561922
rect 75154 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 75774 544350
rect 75154 544226 75774 544294
rect 75154 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 75774 544226
rect 75154 544102 75774 544170
rect 75154 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 75774 544102
rect 75154 543978 75774 544046
rect 75154 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 75774 543978
rect 75154 526350 75774 543922
rect 75154 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 75774 526350
rect 75154 526226 75774 526294
rect 75154 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 75774 526226
rect 75154 526102 75774 526170
rect 75154 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 75774 526102
rect 75154 525978 75774 526046
rect 75154 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 75774 525978
rect 75154 520886 75774 525922
rect 78874 598172 79494 598268
rect 78874 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 79494 598172
rect 78874 598048 79494 598116
rect 78874 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 79494 598048
rect 78874 597924 79494 597992
rect 78874 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 79494 597924
rect 78874 597800 79494 597868
rect 78874 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 79494 597800
rect 78874 586350 79494 597744
rect 78874 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 79494 586350
rect 78874 586226 79494 586294
rect 78874 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 79494 586226
rect 78874 586102 79494 586170
rect 78874 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 79494 586102
rect 78874 585978 79494 586046
rect 78874 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 79494 585978
rect 78874 568350 79494 585922
rect 78874 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 79494 568350
rect 78874 568226 79494 568294
rect 78874 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 79494 568226
rect 78874 568102 79494 568170
rect 78874 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 79494 568102
rect 78874 567978 79494 568046
rect 78874 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 79494 567978
rect 78874 550350 79494 567922
rect 78874 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 79494 550350
rect 78874 550226 79494 550294
rect 78874 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 79494 550226
rect 78874 550102 79494 550170
rect 78874 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 79494 550102
rect 78874 549978 79494 550046
rect 78874 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 79494 549978
rect 78874 532350 79494 549922
rect 78874 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 79494 532350
rect 78874 532226 79494 532294
rect 78874 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 79494 532226
rect 78874 532102 79494 532170
rect 78874 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 79494 532102
rect 78874 531978 79494 532046
rect 78874 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 79494 531978
rect 78874 520886 79494 531922
rect 93154 597212 93774 598268
rect 93154 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 93774 597212
rect 93154 597088 93774 597156
rect 93154 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 93774 597088
rect 93154 596964 93774 597032
rect 93154 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 93774 596964
rect 93154 596840 93774 596908
rect 93154 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 93774 596840
rect 93154 580350 93774 596784
rect 93154 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 93774 580350
rect 93154 580226 93774 580294
rect 93154 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 93774 580226
rect 93154 580102 93774 580170
rect 93154 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 93774 580102
rect 93154 579978 93774 580046
rect 93154 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 93774 579978
rect 93154 562350 93774 579922
rect 93154 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 93774 562350
rect 93154 562226 93774 562294
rect 93154 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 93774 562226
rect 93154 562102 93774 562170
rect 93154 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 93774 562102
rect 93154 561978 93774 562046
rect 93154 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 93774 561978
rect 93154 544350 93774 561922
rect 93154 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 93774 544350
rect 93154 544226 93774 544294
rect 93154 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 93774 544226
rect 93154 544102 93774 544170
rect 93154 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 93774 544102
rect 93154 543978 93774 544046
rect 93154 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 93774 543978
rect 93154 526350 93774 543922
rect 93154 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 93774 526350
rect 93154 526226 93774 526294
rect 93154 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 93774 526226
rect 93154 526102 93774 526170
rect 93154 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 93774 526102
rect 93154 525978 93774 526046
rect 93154 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 93774 525978
rect 93154 520886 93774 525922
rect 96874 598172 97494 598268
rect 96874 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 97494 598172
rect 96874 598048 97494 598116
rect 96874 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 97494 598048
rect 96874 597924 97494 597992
rect 96874 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 97494 597924
rect 96874 597800 97494 597868
rect 96874 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 97494 597800
rect 96874 586350 97494 597744
rect 96874 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 97494 586350
rect 96874 586226 97494 586294
rect 96874 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 97494 586226
rect 96874 586102 97494 586170
rect 96874 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 97494 586102
rect 96874 585978 97494 586046
rect 96874 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 97494 585978
rect 96874 568350 97494 585922
rect 96874 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 97494 568350
rect 96874 568226 97494 568294
rect 96874 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 97494 568226
rect 96874 568102 97494 568170
rect 96874 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 97494 568102
rect 96874 567978 97494 568046
rect 96874 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 97494 567978
rect 96874 550350 97494 567922
rect 96874 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 97494 550350
rect 96874 550226 97494 550294
rect 96874 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 97494 550226
rect 96874 550102 97494 550170
rect 96874 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 97494 550102
rect 96874 549978 97494 550046
rect 96874 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 97494 549978
rect 96874 532350 97494 549922
rect 96874 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 97494 532350
rect 96874 532226 97494 532294
rect 96874 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 97494 532226
rect 96874 532102 97494 532170
rect 96874 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 97494 532102
rect 96874 531978 97494 532046
rect 96874 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 97494 531978
rect 96874 520886 97494 531922
rect 111154 597212 111774 598268
rect 111154 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 111774 597212
rect 111154 597088 111774 597156
rect 111154 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 111774 597088
rect 111154 596964 111774 597032
rect 111154 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 111774 596964
rect 111154 596840 111774 596908
rect 111154 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 111774 596840
rect 111154 580350 111774 596784
rect 111154 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 111774 580350
rect 111154 580226 111774 580294
rect 111154 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 111774 580226
rect 111154 580102 111774 580170
rect 111154 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 111774 580102
rect 111154 579978 111774 580046
rect 111154 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 111774 579978
rect 111154 562350 111774 579922
rect 111154 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 111774 562350
rect 111154 562226 111774 562294
rect 111154 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 111774 562226
rect 111154 562102 111774 562170
rect 111154 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 111774 562102
rect 111154 561978 111774 562046
rect 111154 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 111774 561978
rect 111154 544350 111774 561922
rect 111154 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 111774 544350
rect 111154 544226 111774 544294
rect 111154 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 111774 544226
rect 111154 544102 111774 544170
rect 111154 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 111774 544102
rect 111154 543978 111774 544046
rect 111154 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 111774 543978
rect 111154 526350 111774 543922
rect 111154 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 111774 526350
rect 111154 526226 111774 526294
rect 111154 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 111774 526226
rect 111154 526102 111774 526170
rect 111154 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 111774 526102
rect 111154 525978 111774 526046
rect 111154 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 111774 525978
rect 111154 520886 111774 525922
rect 114874 598172 115494 598268
rect 114874 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 115494 598172
rect 114874 598048 115494 598116
rect 114874 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 115494 598048
rect 114874 597924 115494 597992
rect 114874 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 115494 597924
rect 114874 597800 115494 597868
rect 114874 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 115494 597800
rect 114874 586350 115494 597744
rect 114874 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 115494 586350
rect 114874 586226 115494 586294
rect 114874 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 115494 586226
rect 114874 586102 115494 586170
rect 114874 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 115494 586102
rect 114874 585978 115494 586046
rect 114874 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 115494 585978
rect 114874 568350 115494 585922
rect 114874 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 115494 568350
rect 114874 568226 115494 568294
rect 114874 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 115494 568226
rect 114874 568102 115494 568170
rect 114874 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 115494 568102
rect 114874 567978 115494 568046
rect 114874 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 115494 567978
rect 114874 550350 115494 567922
rect 114874 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 115494 550350
rect 114874 550226 115494 550294
rect 114874 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 115494 550226
rect 114874 550102 115494 550170
rect 114874 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 115494 550102
rect 114874 549978 115494 550046
rect 114874 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 115494 549978
rect 114874 532350 115494 549922
rect 114874 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 115494 532350
rect 114874 532226 115494 532294
rect 114874 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 115494 532226
rect 114874 532102 115494 532170
rect 114874 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 115494 532102
rect 114874 531978 115494 532046
rect 114874 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 115494 531978
rect 114874 520886 115494 531922
rect 129154 597212 129774 598268
rect 129154 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 129774 597212
rect 129154 597088 129774 597156
rect 129154 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 129774 597088
rect 129154 596964 129774 597032
rect 129154 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 129774 596964
rect 129154 596840 129774 596908
rect 129154 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 129774 596840
rect 129154 580350 129774 596784
rect 129154 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 129774 580350
rect 129154 580226 129774 580294
rect 129154 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 129774 580226
rect 129154 580102 129774 580170
rect 129154 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 129774 580102
rect 129154 579978 129774 580046
rect 129154 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 129774 579978
rect 129154 562350 129774 579922
rect 129154 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 129774 562350
rect 129154 562226 129774 562294
rect 129154 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 129774 562226
rect 129154 562102 129774 562170
rect 129154 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 129774 562102
rect 129154 561978 129774 562046
rect 129154 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 129774 561978
rect 129154 544350 129774 561922
rect 129154 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 129774 544350
rect 129154 544226 129774 544294
rect 129154 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 129774 544226
rect 129154 544102 129774 544170
rect 129154 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 129774 544102
rect 129154 543978 129774 544046
rect 129154 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 129774 543978
rect 129154 526350 129774 543922
rect 129154 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 129774 526350
rect 129154 526226 129774 526294
rect 129154 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 129774 526226
rect 129154 526102 129774 526170
rect 129154 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 129774 526102
rect 129154 525978 129774 526046
rect 129154 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 129774 525978
rect 129154 520886 129774 525922
rect 132874 598172 133494 598268
rect 132874 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 133494 598172
rect 132874 598048 133494 598116
rect 132874 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 133494 598048
rect 132874 597924 133494 597992
rect 132874 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 133494 597924
rect 132874 597800 133494 597868
rect 132874 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 133494 597800
rect 132874 586350 133494 597744
rect 132874 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 133494 586350
rect 132874 586226 133494 586294
rect 132874 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 133494 586226
rect 132874 586102 133494 586170
rect 132874 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 133494 586102
rect 132874 585978 133494 586046
rect 132874 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 133494 585978
rect 132874 568350 133494 585922
rect 132874 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 133494 568350
rect 132874 568226 133494 568294
rect 132874 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 133494 568226
rect 132874 568102 133494 568170
rect 132874 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 133494 568102
rect 132874 567978 133494 568046
rect 132874 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 133494 567978
rect 132874 550350 133494 567922
rect 132874 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 133494 550350
rect 132874 550226 133494 550294
rect 132874 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 133494 550226
rect 132874 550102 133494 550170
rect 132874 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 133494 550102
rect 132874 549978 133494 550046
rect 132874 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 133494 549978
rect 132874 532350 133494 549922
rect 132874 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 133494 532350
rect 132874 532226 133494 532294
rect 132874 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 133494 532226
rect 132874 532102 133494 532170
rect 132874 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 133494 532102
rect 132874 531978 133494 532046
rect 132874 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 133494 531978
rect 132874 520886 133494 531922
rect 147154 597212 147774 598268
rect 147154 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 147774 597212
rect 147154 597088 147774 597156
rect 147154 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 147774 597088
rect 147154 596964 147774 597032
rect 147154 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 147774 596964
rect 147154 596840 147774 596908
rect 147154 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 147774 596840
rect 147154 580350 147774 596784
rect 147154 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 147774 580350
rect 147154 580226 147774 580294
rect 147154 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 147774 580226
rect 147154 580102 147774 580170
rect 147154 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 147774 580102
rect 147154 579978 147774 580046
rect 147154 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 147774 579978
rect 147154 562350 147774 579922
rect 147154 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 147774 562350
rect 147154 562226 147774 562294
rect 147154 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 147774 562226
rect 147154 562102 147774 562170
rect 147154 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 147774 562102
rect 147154 561978 147774 562046
rect 147154 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 147774 561978
rect 147154 544350 147774 561922
rect 147154 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 147774 544350
rect 147154 544226 147774 544294
rect 147154 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 147774 544226
rect 147154 544102 147774 544170
rect 147154 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 147774 544102
rect 147154 543978 147774 544046
rect 147154 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 147774 543978
rect 147154 526350 147774 543922
rect 147154 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 147774 526350
rect 147154 526226 147774 526294
rect 147154 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 147774 526226
rect 147154 526102 147774 526170
rect 147154 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 147774 526102
rect 147154 525978 147774 526046
rect 147154 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 147774 525978
rect 147154 520886 147774 525922
rect 150874 598172 151494 598268
rect 150874 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 151494 598172
rect 150874 598048 151494 598116
rect 150874 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 151494 598048
rect 150874 597924 151494 597992
rect 150874 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 151494 597924
rect 150874 597800 151494 597868
rect 150874 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 151494 597800
rect 150874 586350 151494 597744
rect 150874 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 151494 586350
rect 150874 586226 151494 586294
rect 150874 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 151494 586226
rect 150874 586102 151494 586170
rect 150874 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 151494 586102
rect 150874 585978 151494 586046
rect 150874 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 151494 585978
rect 150874 568350 151494 585922
rect 150874 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 151494 568350
rect 150874 568226 151494 568294
rect 150874 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 151494 568226
rect 150874 568102 151494 568170
rect 150874 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 151494 568102
rect 150874 567978 151494 568046
rect 150874 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 151494 567978
rect 150874 550350 151494 567922
rect 150874 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 151494 550350
rect 150874 550226 151494 550294
rect 150874 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 151494 550226
rect 150874 550102 151494 550170
rect 150874 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 151494 550102
rect 150874 549978 151494 550046
rect 150874 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 151494 549978
rect 150874 532350 151494 549922
rect 150874 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 151494 532350
rect 150874 532226 151494 532294
rect 150874 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 151494 532226
rect 150874 532102 151494 532170
rect 150874 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 151494 532102
rect 150874 531978 151494 532046
rect 150874 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 151494 531978
rect 150874 520886 151494 531922
rect 165154 597212 165774 598268
rect 165154 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 165774 597212
rect 165154 597088 165774 597156
rect 165154 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 165774 597088
rect 165154 596964 165774 597032
rect 165154 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 165774 596964
rect 165154 596840 165774 596908
rect 165154 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 165774 596840
rect 165154 580350 165774 596784
rect 165154 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 165774 580350
rect 165154 580226 165774 580294
rect 165154 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 165774 580226
rect 165154 580102 165774 580170
rect 165154 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 165774 580102
rect 165154 579978 165774 580046
rect 165154 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 165774 579978
rect 165154 562350 165774 579922
rect 165154 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 165774 562350
rect 165154 562226 165774 562294
rect 165154 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 165774 562226
rect 165154 562102 165774 562170
rect 165154 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 165774 562102
rect 165154 561978 165774 562046
rect 165154 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 165774 561978
rect 165154 544350 165774 561922
rect 165154 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 165774 544350
rect 165154 544226 165774 544294
rect 165154 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 165774 544226
rect 165154 544102 165774 544170
rect 165154 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 165774 544102
rect 165154 543978 165774 544046
rect 165154 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 165774 543978
rect 165154 526350 165774 543922
rect 165154 526294 165250 526350
rect 165306 526294 165374 526350
rect 165430 526294 165498 526350
rect 165554 526294 165622 526350
rect 165678 526294 165774 526350
rect 165154 526226 165774 526294
rect 165154 526170 165250 526226
rect 165306 526170 165374 526226
rect 165430 526170 165498 526226
rect 165554 526170 165622 526226
rect 165678 526170 165774 526226
rect 165154 526102 165774 526170
rect 165154 526046 165250 526102
rect 165306 526046 165374 526102
rect 165430 526046 165498 526102
rect 165554 526046 165622 526102
rect 165678 526046 165774 526102
rect 165154 525978 165774 526046
rect 165154 525922 165250 525978
rect 165306 525922 165374 525978
rect 165430 525922 165498 525978
rect 165554 525922 165622 525978
rect 165678 525922 165774 525978
rect 165154 520886 165774 525922
rect 168874 598172 169494 598268
rect 168874 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 169494 598172
rect 168874 598048 169494 598116
rect 168874 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 169494 598048
rect 168874 597924 169494 597992
rect 168874 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 169494 597924
rect 168874 597800 169494 597868
rect 168874 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 169494 597800
rect 168874 586350 169494 597744
rect 168874 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 169494 586350
rect 168874 586226 169494 586294
rect 168874 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 169494 586226
rect 168874 586102 169494 586170
rect 168874 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 169494 586102
rect 168874 585978 169494 586046
rect 168874 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 169494 585978
rect 168874 568350 169494 585922
rect 168874 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 169494 568350
rect 168874 568226 169494 568294
rect 168874 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 169494 568226
rect 168874 568102 169494 568170
rect 168874 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 169494 568102
rect 168874 567978 169494 568046
rect 168874 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 169494 567978
rect 168874 550350 169494 567922
rect 168874 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 169494 550350
rect 168874 550226 169494 550294
rect 168874 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 169494 550226
rect 168874 550102 169494 550170
rect 168874 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 169494 550102
rect 168874 549978 169494 550046
rect 168874 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 169494 549978
rect 168874 532350 169494 549922
rect 168874 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 169494 532350
rect 168874 532226 169494 532294
rect 168874 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 169494 532226
rect 168874 532102 169494 532170
rect 168874 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 169494 532102
rect 168874 531978 169494 532046
rect 168874 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 169494 531978
rect 168874 520886 169494 531922
rect 183154 597212 183774 598268
rect 183154 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 183774 597212
rect 183154 597088 183774 597156
rect 183154 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 183774 597088
rect 183154 596964 183774 597032
rect 183154 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 183774 596964
rect 183154 596840 183774 596908
rect 183154 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 183774 596840
rect 183154 580350 183774 596784
rect 183154 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 183774 580350
rect 183154 580226 183774 580294
rect 183154 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 183774 580226
rect 183154 580102 183774 580170
rect 183154 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 183774 580102
rect 183154 579978 183774 580046
rect 183154 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 183774 579978
rect 183154 562350 183774 579922
rect 183154 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 183774 562350
rect 183154 562226 183774 562294
rect 183154 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 183774 562226
rect 183154 562102 183774 562170
rect 183154 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 183774 562102
rect 183154 561978 183774 562046
rect 183154 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 183774 561978
rect 183154 544350 183774 561922
rect 183154 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 183774 544350
rect 183154 544226 183774 544294
rect 183154 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 183774 544226
rect 183154 544102 183774 544170
rect 183154 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 183774 544102
rect 183154 543978 183774 544046
rect 183154 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 183774 543978
rect 183154 526350 183774 543922
rect 183154 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 183774 526350
rect 183154 526226 183774 526294
rect 183154 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 183774 526226
rect 183154 526102 183774 526170
rect 183154 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 183774 526102
rect 183154 525978 183774 526046
rect 183154 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 183774 525978
rect 183154 520886 183774 525922
rect 186874 598172 187494 598268
rect 186874 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 187494 598172
rect 186874 598048 187494 598116
rect 186874 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 187494 598048
rect 186874 597924 187494 597992
rect 186874 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 187494 597924
rect 186874 597800 187494 597868
rect 186874 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 187494 597800
rect 186874 586350 187494 597744
rect 186874 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 187494 586350
rect 186874 586226 187494 586294
rect 186874 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 187494 586226
rect 186874 586102 187494 586170
rect 186874 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 187494 586102
rect 186874 585978 187494 586046
rect 186874 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 187494 585978
rect 186874 568350 187494 585922
rect 186874 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 187494 568350
rect 186874 568226 187494 568294
rect 186874 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 187494 568226
rect 186874 568102 187494 568170
rect 186874 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 187494 568102
rect 186874 567978 187494 568046
rect 186874 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 187494 567978
rect 186874 550350 187494 567922
rect 186874 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 187494 550350
rect 186874 550226 187494 550294
rect 186874 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 187494 550226
rect 186874 550102 187494 550170
rect 186874 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 187494 550102
rect 186874 549978 187494 550046
rect 186874 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 187494 549978
rect 186874 532350 187494 549922
rect 186874 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 187494 532350
rect 186874 532226 187494 532294
rect 186874 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 187494 532226
rect 186874 532102 187494 532170
rect 186874 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 187494 532102
rect 186874 531978 187494 532046
rect 186874 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 187494 531978
rect 186874 520886 187494 531922
rect 201154 597212 201774 598268
rect 201154 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 201774 597212
rect 201154 597088 201774 597156
rect 201154 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 201774 597088
rect 201154 596964 201774 597032
rect 201154 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 201774 596964
rect 201154 596840 201774 596908
rect 201154 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 201774 596840
rect 201154 580350 201774 596784
rect 201154 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 201774 580350
rect 201154 580226 201774 580294
rect 201154 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 201774 580226
rect 201154 580102 201774 580170
rect 201154 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 201774 580102
rect 201154 579978 201774 580046
rect 201154 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 201774 579978
rect 201154 562350 201774 579922
rect 201154 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 201774 562350
rect 201154 562226 201774 562294
rect 201154 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 201774 562226
rect 201154 562102 201774 562170
rect 201154 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 201774 562102
rect 201154 561978 201774 562046
rect 201154 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 201774 561978
rect 201154 544350 201774 561922
rect 201154 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 201774 544350
rect 201154 544226 201774 544294
rect 201154 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 201774 544226
rect 201154 544102 201774 544170
rect 201154 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 201774 544102
rect 201154 543978 201774 544046
rect 201154 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 201774 543978
rect 201154 526350 201774 543922
rect 201154 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 201774 526350
rect 201154 526226 201774 526294
rect 201154 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 201774 526226
rect 201154 526102 201774 526170
rect 201154 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 201774 526102
rect 201154 525978 201774 526046
rect 201154 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 201774 525978
rect 201154 520886 201774 525922
rect 204874 598172 205494 598268
rect 204874 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 205494 598172
rect 204874 598048 205494 598116
rect 204874 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 205494 598048
rect 204874 597924 205494 597992
rect 204874 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 205494 597924
rect 204874 597800 205494 597868
rect 204874 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 205494 597800
rect 204874 586350 205494 597744
rect 204874 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 205494 586350
rect 204874 586226 205494 586294
rect 204874 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 205494 586226
rect 204874 586102 205494 586170
rect 204874 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 205494 586102
rect 204874 585978 205494 586046
rect 204874 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 205494 585978
rect 204874 568350 205494 585922
rect 204874 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 205494 568350
rect 204874 568226 205494 568294
rect 204874 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 205494 568226
rect 204874 568102 205494 568170
rect 204874 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 205494 568102
rect 204874 567978 205494 568046
rect 204874 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 205494 567978
rect 204874 550350 205494 567922
rect 204874 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 205494 550350
rect 204874 550226 205494 550294
rect 204874 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 205494 550226
rect 204874 550102 205494 550170
rect 204874 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 205494 550102
rect 204874 549978 205494 550046
rect 204874 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 205494 549978
rect 204874 532350 205494 549922
rect 204874 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 205494 532350
rect 204874 532226 205494 532294
rect 204874 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 205494 532226
rect 204874 532102 205494 532170
rect 204874 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 205494 532102
rect 204874 531978 205494 532046
rect 204874 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 205494 531978
rect 204874 520886 205494 531922
rect 219154 597212 219774 598268
rect 219154 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 219774 597212
rect 219154 597088 219774 597156
rect 219154 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 219774 597088
rect 219154 596964 219774 597032
rect 219154 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 219774 596964
rect 219154 596840 219774 596908
rect 219154 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 219774 596840
rect 219154 580350 219774 596784
rect 219154 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 219774 580350
rect 219154 580226 219774 580294
rect 219154 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 219774 580226
rect 219154 580102 219774 580170
rect 219154 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 219774 580102
rect 219154 579978 219774 580046
rect 219154 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 219774 579978
rect 219154 562350 219774 579922
rect 219154 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 219774 562350
rect 219154 562226 219774 562294
rect 219154 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 219774 562226
rect 219154 562102 219774 562170
rect 219154 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 219774 562102
rect 219154 561978 219774 562046
rect 219154 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 219774 561978
rect 219154 544350 219774 561922
rect 219154 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 219774 544350
rect 219154 544226 219774 544294
rect 219154 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 219774 544226
rect 219154 544102 219774 544170
rect 219154 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 219774 544102
rect 219154 543978 219774 544046
rect 219154 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 219774 543978
rect 219154 526350 219774 543922
rect 219154 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 219774 526350
rect 219154 526226 219774 526294
rect 219154 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 219774 526226
rect 219154 526102 219774 526170
rect 219154 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 219774 526102
rect 219154 525978 219774 526046
rect 219154 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 219774 525978
rect 219154 520886 219774 525922
rect 222874 598172 223494 598268
rect 222874 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 223494 598172
rect 222874 598048 223494 598116
rect 222874 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 223494 598048
rect 222874 597924 223494 597992
rect 222874 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 223494 597924
rect 222874 597800 223494 597868
rect 222874 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 223494 597800
rect 222874 586350 223494 597744
rect 222874 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 223494 586350
rect 222874 586226 223494 586294
rect 222874 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 223494 586226
rect 222874 586102 223494 586170
rect 222874 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 223494 586102
rect 222874 585978 223494 586046
rect 222874 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 223494 585978
rect 222874 568350 223494 585922
rect 222874 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 223494 568350
rect 222874 568226 223494 568294
rect 222874 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 223494 568226
rect 222874 568102 223494 568170
rect 222874 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 223494 568102
rect 222874 567978 223494 568046
rect 222874 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 223494 567978
rect 222874 550350 223494 567922
rect 222874 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 223494 550350
rect 222874 550226 223494 550294
rect 222874 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 223494 550226
rect 222874 550102 223494 550170
rect 222874 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 223494 550102
rect 222874 549978 223494 550046
rect 222874 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 223494 549978
rect 222874 532350 223494 549922
rect 222874 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 223494 532350
rect 222874 532226 223494 532294
rect 222874 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 223494 532226
rect 222874 532102 223494 532170
rect 222874 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 223494 532102
rect 222874 531978 223494 532046
rect 222874 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 223494 531978
rect 222874 520886 223494 531922
rect 237154 597212 237774 598268
rect 237154 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 237774 597212
rect 237154 597088 237774 597156
rect 237154 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 237774 597088
rect 237154 596964 237774 597032
rect 237154 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 237774 596964
rect 237154 596840 237774 596908
rect 237154 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 237774 596840
rect 237154 580350 237774 596784
rect 237154 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 237774 580350
rect 237154 580226 237774 580294
rect 237154 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 237774 580226
rect 237154 580102 237774 580170
rect 237154 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 237774 580102
rect 237154 579978 237774 580046
rect 237154 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 237774 579978
rect 237154 562350 237774 579922
rect 237154 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 237774 562350
rect 237154 562226 237774 562294
rect 237154 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 237774 562226
rect 237154 562102 237774 562170
rect 237154 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 237774 562102
rect 237154 561978 237774 562046
rect 237154 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 237774 561978
rect 237154 544350 237774 561922
rect 237154 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 237774 544350
rect 237154 544226 237774 544294
rect 237154 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 237774 544226
rect 237154 544102 237774 544170
rect 237154 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 237774 544102
rect 237154 543978 237774 544046
rect 237154 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 237774 543978
rect 237154 526350 237774 543922
rect 237154 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 237774 526350
rect 237154 526226 237774 526294
rect 237154 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 237774 526226
rect 237154 526102 237774 526170
rect 237154 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 237774 526102
rect 237154 525978 237774 526046
rect 237154 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 237774 525978
rect 237154 520886 237774 525922
rect 240874 598172 241494 598268
rect 240874 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 241494 598172
rect 240874 598048 241494 598116
rect 240874 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 241494 598048
rect 240874 597924 241494 597992
rect 240874 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 241494 597924
rect 240874 597800 241494 597868
rect 240874 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 241494 597800
rect 240874 586350 241494 597744
rect 240874 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 241494 586350
rect 240874 586226 241494 586294
rect 240874 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 241494 586226
rect 240874 586102 241494 586170
rect 240874 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 241494 586102
rect 240874 585978 241494 586046
rect 240874 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 241494 585978
rect 240874 568350 241494 585922
rect 240874 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 241494 568350
rect 240874 568226 241494 568294
rect 240874 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 241494 568226
rect 240874 568102 241494 568170
rect 240874 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 241494 568102
rect 240874 567978 241494 568046
rect 240874 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 241494 567978
rect 240874 550350 241494 567922
rect 240874 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 241494 550350
rect 240874 550226 241494 550294
rect 240874 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 241494 550226
rect 240874 550102 241494 550170
rect 240874 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 241494 550102
rect 240874 549978 241494 550046
rect 240874 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 241494 549978
rect 240874 532350 241494 549922
rect 240874 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 241494 532350
rect 240874 532226 241494 532294
rect 240874 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 241494 532226
rect 240874 532102 241494 532170
rect 240874 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 241494 532102
rect 240874 531978 241494 532046
rect 240874 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 241494 531978
rect 240874 520886 241494 531922
rect 255154 597212 255774 598268
rect 255154 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 255774 597212
rect 255154 597088 255774 597156
rect 255154 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 255774 597088
rect 255154 596964 255774 597032
rect 255154 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 255774 596964
rect 255154 596840 255774 596908
rect 255154 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 255774 596840
rect 255154 580350 255774 596784
rect 255154 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 255774 580350
rect 255154 580226 255774 580294
rect 255154 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 255774 580226
rect 255154 580102 255774 580170
rect 255154 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 255774 580102
rect 255154 579978 255774 580046
rect 255154 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 255774 579978
rect 255154 562350 255774 579922
rect 255154 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 255774 562350
rect 255154 562226 255774 562294
rect 255154 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 255774 562226
rect 255154 562102 255774 562170
rect 255154 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 255774 562102
rect 255154 561978 255774 562046
rect 255154 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 255774 561978
rect 255154 544350 255774 561922
rect 255154 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 255774 544350
rect 255154 544226 255774 544294
rect 255154 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 255774 544226
rect 255154 544102 255774 544170
rect 255154 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 255774 544102
rect 255154 543978 255774 544046
rect 255154 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 255774 543978
rect 255154 526350 255774 543922
rect 255154 526294 255250 526350
rect 255306 526294 255374 526350
rect 255430 526294 255498 526350
rect 255554 526294 255622 526350
rect 255678 526294 255774 526350
rect 255154 526226 255774 526294
rect 255154 526170 255250 526226
rect 255306 526170 255374 526226
rect 255430 526170 255498 526226
rect 255554 526170 255622 526226
rect 255678 526170 255774 526226
rect 255154 526102 255774 526170
rect 255154 526046 255250 526102
rect 255306 526046 255374 526102
rect 255430 526046 255498 526102
rect 255554 526046 255622 526102
rect 255678 526046 255774 526102
rect 255154 525978 255774 526046
rect 255154 525922 255250 525978
rect 255306 525922 255374 525978
rect 255430 525922 255498 525978
rect 255554 525922 255622 525978
rect 255678 525922 255774 525978
rect 255154 520886 255774 525922
rect 258874 598172 259494 598268
rect 258874 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 259494 598172
rect 258874 598048 259494 598116
rect 258874 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 259494 598048
rect 258874 597924 259494 597992
rect 258874 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 259494 597924
rect 258874 597800 259494 597868
rect 258874 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 259494 597800
rect 258874 586350 259494 597744
rect 258874 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 259494 586350
rect 258874 586226 259494 586294
rect 258874 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 259494 586226
rect 258874 586102 259494 586170
rect 258874 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 259494 586102
rect 258874 585978 259494 586046
rect 258874 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 259494 585978
rect 258874 568350 259494 585922
rect 258874 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 259494 568350
rect 258874 568226 259494 568294
rect 258874 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 259494 568226
rect 258874 568102 259494 568170
rect 258874 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 259494 568102
rect 258874 567978 259494 568046
rect 258874 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 259494 567978
rect 258874 550350 259494 567922
rect 258874 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 259494 550350
rect 258874 550226 259494 550294
rect 258874 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 259494 550226
rect 258874 550102 259494 550170
rect 258874 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 259494 550102
rect 258874 549978 259494 550046
rect 258874 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 259494 549978
rect 258874 532350 259494 549922
rect 258874 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 259494 532350
rect 258874 532226 259494 532294
rect 258874 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 259494 532226
rect 258874 532102 259494 532170
rect 258874 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 259494 532102
rect 258874 531978 259494 532046
rect 258874 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 259494 531978
rect 258874 520886 259494 531922
rect 273154 597212 273774 598268
rect 273154 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 273774 597212
rect 273154 597088 273774 597156
rect 273154 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 273774 597088
rect 273154 596964 273774 597032
rect 273154 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 273774 596964
rect 273154 596840 273774 596908
rect 273154 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 273774 596840
rect 273154 580350 273774 596784
rect 273154 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 273774 580350
rect 273154 580226 273774 580294
rect 273154 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 273774 580226
rect 273154 580102 273774 580170
rect 273154 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 273774 580102
rect 273154 579978 273774 580046
rect 273154 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 273774 579978
rect 273154 562350 273774 579922
rect 273154 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 273774 562350
rect 273154 562226 273774 562294
rect 273154 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 273774 562226
rect 273154 562102 273774 562170
rect 273154 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 273774 562102
rect 273154 561978 273774 562046
rect 273154 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 273774 561978
rect 273154 544350 273774 561922
rect 273154 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 273774 544350
rect 273154 544226 273774 544294
rect 273154 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 273774 544226
rect 273154 544102 273774 544170
rect 273154 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 273774 544102
rect 273154 543978 273774 544046
rect 273154 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 273774 543978
rect 273154 526350 273774 543922
rect 273154 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 273774 526350
rect 273154 526226 273774 526294
rect 273154 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 273774 526226
rect 273154 526102 273774 526170
rect 273154 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 273774 526102
rect 273154 525978 273774 526046
rect 273154 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 273774 525978
rect 273154 520886 273774 525922
rect 276874 598172 277494 598268
rect 276874 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 277494 598172
rect 276874 598048 277494 598116
rect 276874 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 277494 598048
rect 276874 597924 277494 597992
rect 276874 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 277494 597924
rect 276874 597800 277494 597868
rect 276874 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 277494 597800
rect 276874 586350 277494 597744
rect 276874 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 277494 586350
rect 276874 586226 277494 586294
rect 276874 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 277494 586226
rect 276874 586102 277494 586170
rect 276874 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 277494 586102
rect 276874 585978 277494 586046
rect 276874 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 277494 585978
rect 276874 568350 277494 585922
rect 276874 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 277494 568350
rect 276874 568226 277494 568294
rect 276874 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 277494 568226
rect 276874 568102 277494 568170
rect 276874 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 277494 568102
rect 276874 567978 277494 568046
rect 276874 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 277494 567978
rect 276874 550350 277494 567922
rect 276874 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 277494 550350
rect 276874 550226 277494 550294
rect 276874 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 277494 550226
rect 276874 550102 277494 550170
rect 276874 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 277494 550102
rect 276874 549978 277494 550046
rect 276874 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 277494 549978
rect 276874 532350 277494 549922
rect 276874 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 277494 532350
rect 276874 532226 277494 532294
rect 276874 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 277494 532226
rect 276874 532102 277494 532170
rect 276874 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 277494 532102
rect 276874 531978 277494 532046
rect 276874 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 277494 531978
rect 276874 520886 277494 531922
rect 291154 597212 291774 598268
rect 291154 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 291774 597212
rect 291154 597088 291774 597156
rect 291154 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 291774 597088
rect 291154 596964 291774 597032
rect 291154 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 291774 596964
rect 291154 596840 291774 596908
rect 291154 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 291774 596840
rect 291154 580350 291774 596784
rect 291154 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 291774 580350
rect 291154 580226 291774 580294
rect 291154 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 291774 580226
rect 291154 580102 291774 580170
rect 291154 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 291774 580102
rect 291154 579978 291774 580046
rect 291154 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 291774 579978
rect 291154 562350 291774 579922
rect 291154 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 291774 562350
rect 291154 562226 291774 562294
rect 291154 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 291774 562226
rect 291154 562102 291774 562170
rect 291154 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 291774 562102
rect 291154 561978 291774 562046
rect 291154 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 291774 561978
rect 291154 544350 291774 561922
rect 291154 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 291774 544350
rect 291154 544226 291774 544294
rect 291154 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 291774 544226
rect 291154 544102 291774 544170
rect 291154 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 291774 544102
rect 291154 543978 291774 544046
rect 291154 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 291774 543978
rect 291154 526350 291774 543922
rect 291154 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 291774 526350
rect 291154 526226 291774 526294
rect 291154 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 291774 526226
rect 291154 526102 291774 526170
rect 291154 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 291774 526102
rect 291154 525978 291774 526046
rect 291154 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 291774 525978
rect 291154 520886 291774 525922
rect 294874 598172 295494 598268
rect 294874 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 295494 598172
rect 294874 598048 295494 598116
rect 294874 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 295494 598048
rect 294874 597924 295494 597992
rect 294874 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 295494 597924
rect 294874 597800 295494 597868
rect 294874 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 295494 597800
rect 294874 586350 295494 597744
rect 294874 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 295494 586350
rect 294874 586226 295494 586294
rect 294874 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 295494 586226
rect 294874 586102 295494 586170
rect 294874 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 295494 586102
rect 294874 585978 295494 586046
rect 294874 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 295494 585978
rect 294874 568350 295494 585922
rect 294874 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 295494 568350
rect 294874 568226 295494 568294
rect 294874 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 295494 568226
rect 294874 568102 295494 568170
rect 294874 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 295494 568102
rect 294874 567978 295494 568046
rect 294874 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 295494 567978
rect 294874 550350 295494 567922
rect 294874 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 295494 550350
rect 294874 550226 295494 550294
rect 294874 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 295494 550226
rect 294874 550102 295494 550170
rect 294874 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 295494 550102
rect 294874 549978 295494 550046
rect 294874 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 295494 549978
rect 294874 532350 295494 549922
rect 294874 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 295494 532350
rect 294874 532226 295494 532294
rect 294874 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 295494 532226
rect 294874 532102 295494 532170
rect 294874 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 295494 532102
rect 294874 531978 295494 532046
rect 294874 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 295494 531978
rect 294874 520886 295494 531922
rect 309154 597212 309774 598268
rect 309154 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 309774 597212
rect 309154 597088 309774 597156
rect 309154 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 309774 597088
rect 309154 596964 309774 597032
rect 309154 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 309774 596964
rect 309154 596840 309774 596908
rect 309154 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 309774 596840
rect 309154 580350 309774 596784
rect 309154 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 309774 580350
rect 309154 580226 309774 580294
rect 309154 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 309774 580226
rect 309154 580102 309774 580170
rect 309154 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 309774 580102
rect 309154 579978 309774 580046
rect 309154 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 309774 579978
rect 309154 562350 309774 579922
rect 309154 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 309774 562350
rect 309154 562226 309774 562294
rect 309154 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 309774 562226
rect 309154 562102 309774 562170
rect 309154 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 309774 562102
rect 309154 561978 309774 562046
rect 309154 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 309774 561978
rect 309154 544350 309774 561922
rect 309154 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 309774 544350
rect 309154 544226 309774 544294
rect 309154 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 309774 544226
rect 309154 544102 309774 544170
rect 309154 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 309774 544102
rect 309154 543978 309774 544046
rect 309154 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 309774 543978
rect 309154 526350 309774 543922
rect 309154 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 309774 526350
rect 309154 526226 309774 526294
rect 309154 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 309774 526226
rect 309154 526102 309774 526170
rect 309154 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 309774 526102
rect 309154 525978 309774 526046
rect 309154 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 309774 525978
rect 309154 520886 309774 525922
rect 312874 598172 313494 598268
rect 312874 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 313494 598172
rect 312874 598048 313494 598116
rect 312874 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 313494 598048
rect 312874 597924 313494 597992
rect 312874 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 313494 597924
rect 312874 597800 313494 597868
rect 312874 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 313494 597800
rect 312874 586350 313494 597744
rect 312874 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 313494 586350
rect 312874 586226 313494 586294
rect 312874 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 313494 586226
rect 312874 586102 313494 586170
rect 312874 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 313494 586102
rect 312874 585978 313494 586046
rect 312874 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 313494 585978
rect 312874 568350 313494 585922
rect 312874 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 313494 568350
rect 312874 568226 313494 568294
rect 312874 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 313494 568226
rect 312874 568102 313494 568170
rect 312874 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 313494 568102
rect 312874 567978 313494 568046
rect 312874 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 313494 567978
rect 312874 550350 313494 567922
rect 312874 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 313494 550350
rect 312874 550226 313494 550294
rect 312874 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 313494 550226
rect 312874 550102 313494 550170
rect 312874 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 313494 550102
rect 312874 549978 313494 550046
rect 312874 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 313494 549978
rect 312874 532350 313494 549922
rect 312874 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 313494 532350
rect 312874 532226 313494 532294
rect 312874 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 313494 532226
rect 312874 532102 313494 532170
rect 312874 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 313494 532102
rect 312874 531978 313494 532046
rect 312874 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 313494 531978
rect 312874 520886 313494 531922
rect 327154 597212 327774 598268
rect 327154 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 327774 597212
rect 327154 597088 327774 597156
rect 327154 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 327774 597088
rect 327154 596964 327774 597032
rect 327154 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 327774 596964
rect 327154 596840 327774 596908
rect 327154 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 327774 596840
rect 327154 580350 327774 596784
rect 327154 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 327774 580350
rect 327154 580226 327774 580294
rect 327154 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 327774 580226
rect 327154 580102 327774 580170
rect 327154 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 327774 580102
rect 327154 579978 327774 580046
rect 327154 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 327774 579978
rect 327154 562350 327774 579922
rect 327154 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 327774 562350
rect 327154 562226 327774 562294
rect 327154 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 327774 562226
rect 327154 562102 327774 562170
rect 327154 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 327774 562102
rect 327154 561978 327774 562046
rect 327154 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 327774 561978
rect 327154 544350 327774 561922
rect 327154 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 327774 544350
rect 327154 544226 327774 544294
rect 327154 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 327774 544226
rect 327154 544102 327774 544170
rect 327154 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 327774 544102
rect 327154 543978 327774 544046
rect 327154 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 327774 543978
rect 327154 526350 327774 543922
rect 327154 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 327774 526350
rect 327154 526226 327774 526294
rect 327154 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 327774 526226
rect 327154 526102 327774 526170
rect 327154 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 327774 526102
rect 327154 525978 327774 526046
rect 327154 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 327774 525978
rect 327154 520886 327774 525922
rect 330874 598172 331494 598268
rect 330874 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 331494 598172
rect 330874 598048 331494 598116
rect 330874 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 331494 598048
rect 330874 597924 331494 597992
rect 330874 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 331494 597924
rect 330874 597800 331494 597868
rect 330874 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 331494 597800
rect 330874 586350 331494 597744
rect 330874 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 331494 586350
rect 330874 586226 331494 586294
rect 330874 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 331494 586226
rect 330874 586102 331494 586170
rect 330874 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 331494 586102
rect 330874 585978 331494 586046
rect 330874 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 331494 585978
rect 330874 568350 331494 585922
rect 330874 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 331494 568350
rect 330874 568226 331494 568294
rect 330874 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 331494 568226
rect 330874 568102 331494 568170
rect 330874 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 331494 568102
rect 330874 567978 331494 568046
rect 330874 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 331494 567978
rect 330874 550350 331494 567922
rect 330874 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 331494 550350
rect 330874 550226 331494 550294
rect 330874 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 331494 550226
rect 330874 550102 331494 550170
rect 330874 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 331494 550102
rect 330874 549978 331494 550046
rect 330874 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 331494 549978
rect 330874 532350 331494 549922
rect 330874 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 331494 532350
rect 330874 532226 331494 532294
rect 330874 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 331494 532226
rect 330874 532102 331494 532170
rect 330874 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 331494 532102
rect 330874 531978 331494 532046
rect 330874 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 331494 531978
rect 330874 520886 331494 531922
rect 345154 597212 345774 598268
rect 345154 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 345774 597212
rect 345154 597088 345774 597156
rect 345154 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 345774 597088
rect 345154 596964 345774 597032
rect 345154 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 345774 596964
rect 345154 596840 345774 596908
rect 345154 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 345774 596840
rect 345154 580350 345774 596784
rect 345154 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 345774 580350
rect 345154 580226 345774 580294
rect 345154 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 345774 580226
rect 345154 580102 345774 580170
rect 345154 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 345774 580102
rect 345154 579978 345774 580046
rect 345154 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 345774 579978
rect 345154 562350 345774 579922
rect 345154 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 345774 562350
rect 345154 562226 345774 562294
rect 345154 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 345774 562226
rect 345154 562102 345774 562170
rect 345154 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 345774 562102
rect 345154 561978 345774 562046
rect 345154 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 345774 561978
rect 345154 544350 345774 561922
rect 345154 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 345774 544350
rect 345154 544226 345774 544294
rect 345154 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 345774 544226
rect 345154 544102 345774 544170
rect 345154 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 345774 544102
rect 345154 543978 345774 544046
rect 345154 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 345774 543978
rect 345154 526350 345774 543922
rect 345154 526294 345250 526350
rect 345306 526294 345374 526350
rect 345430 526294 345498 526350
rect 345554 526294 345622 526350
rect 345678 526294 345774 526350
rect 345154 526226 345774 526294
rect 345154 526170 345250 526226
rect 345306 526170 345374 526226
rect 345430 526170 345498 526226
rect 345554 526170 345622 526226
rect 345678 526170 345774 526226
rect 345154 526102 345774 526170
rect 345154 526046 345250 526102
rect 345306 526046 345374 526102
rect 345430 526046 345498 526102
rect 345554 526046 345622 526102
rect 345678 526046 345774 526102
rect 345154 525978 345774 526046
rect 345154 525922 345250 525978
rect 345306 525922 345374 525978
rect 345430 525922 345498 525978
rect 345554 525922 345622 525978
rect 345678 525922 345774 525978
rect 345154 520886 345774 525922
rect 348874 598172 349494 598268
rect 348874 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 349494 598172
rect 348874 598048 349494 598116
rect 348874 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 349494 598048
rect 348874 597924 349494 597992
rect 348874 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 349494 597924
rect 348874 597800 349494 597868
rect 348874 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 349494 597800
rect 348874 586350 349494 597744
rect 348874 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 349494 586350
rect 348874 586226 349494 586294
rect 348874 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 349494 586226
rect 348874 586102 349494 586170
rect 348874 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 349494 586102
rect 348874 585978 349494 586046
rect 348874 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 349494 585978
rect 348874 568350 349494 585922
rect 348874 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 349494 568350
rect 348874 568226 349494 568294
rect 348874 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 349494 568226
rect 348874 568102 349494 568170
rect 348874 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 349494 568102
rect 348874 567978 349494 568046
rect 348874 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 349494 567978
rect 348874 550350 349494 567922
rect 348874 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 349494 550350
rect 348874 550226 349494 550294
rect 348874 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 349494 550226
rect 348874 550102 349494 550170
rect 348874 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 349494 550102
rect 348874 549978 349494 550046
rect 348874 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 349494 549978
rect 348874 532350 349494 549922
rect 348874 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 349494 532350
rect 348874 532226 349494 532294
rect 348874 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 349494 532226
rect 348874 532102 349494 532170
rect 348874 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 349494 532102
rect 348874 531978 349494 532046
rect 348874 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 349494 531978
rect 348874 520886 349494 531922
rect 363154 597212 363774 598268
rect 363154 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 363774 597212
rect 363154 597088 363774 597156
rect 363154 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 363774 597088
rect 363154 596964 363774 597032
rect 363154 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 363774 596964
rect 363154 596840 363774 596908
rect 363154 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 363774 596840
rect 363154 580350 363774 596784
rect 363154 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 363774 580350
rect 363154 580226 363774 580294
rect 363154 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 363774 580226
rect 363154 580102 363774 580170
rect 363154 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 363774 580102
rect 363154 579978 363774 580046
rect 363154 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 363774 579978
rect 363154 562350 363774 579922
rect 363154 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 363774 562350
rect 363154 562226 363774 562294
rect 363154 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 363774 562226
rect 363154 562102 363774 562170
rect 363154 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 363774 562102
rect 363154 561978 363774 562046
rect 363154 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 363774 561978
rect 363154 544350 363774 561922
rect 363154 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 363774 544350
rect 363154 544226 363774 544294
rect 363154 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 363774 544226
rect 363154 544102 363774 544170
rect 363154 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 363774 544102
rect 363154 543978 363774 544046
rect 363154 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 363774 543978
rect 363154 526350 363774 543922
rect 363154 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 363774 526350
rect 363154 526226 363774 526294
rect 363154 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 363774 526226
rect 363154 526102 363774 526170
rect 363154 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 363774 526102
rect 363154 525978 363774 526046
rect 363154 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 363774 525978
rect 363154 520886 363774 525922
rect 366874 598172 367494 598268
rect 366874 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 367494 598172
rect 366874 598048 367494 598116
rect 366874 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 367494 598048
rect 366874 597924 367494 597992
rect 366874 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 367494 597924
rect 366874 597800 367494 597868
rect 366874 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 367494 597800
rect 366874 586350 367494 597744
rect 366874 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 367494 586350
rect 366874 586226 367494 586294
rect 366874 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 367494 586226
rect 366874 586102 367494 586170
rect 366874 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 367494 586102
rect 366874 585978 367494 586046
rect 366874 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 367494 585978
rect 366874 568350 367494 585922
rect 366874 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 367494 568350
rect 366874 568226 367494 568294
rect 366874 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 367494 568226
rect 366874 568102 367494 568170
rect 366874 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 367494 568102
rect 366874 567978 367494 568046
rect 366874 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 367494 567978
rect 366874 550350 367494 567922
rect 366874 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 367494 550350
rect 366874 550226 367494 550294
rect 366874 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 367494 550226
rect 366874 550102 367494 550170
rect 366874 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 367494 550102
rect 366874 549978 367494 550046
rect 366874 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 367494 549978
rect 366874 532350 367494 549922
rect 366874 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 367494 532350
rect 366874 532226 367494 532294
rect 366874 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 367494 532226
rect 366874 532102 367494 532170
rect 366874 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 367494 532102
rect 366874 531978 367494 532046
rect 366874 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 367494 531978
rect 366874 520886 367494 531922
rect 381154 597212 381774 598268
rect 381154 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 381774 597212
rect 381154 597088 381774 597156
rect 381154 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 381774 597088
rect 381154 596964 381774 597032
rect 381154 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 381774 596964
rect 381154 596840 381774 596908
rect 381154 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 381774 596840
rect 381154 580350 381774 596784
rect 381154 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 381774 580350
rect 381154 580226 381774 580294
rect 381154 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 381774 580226
rect 381154 580102 381774 580170
rect 381154 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 381774 580102
rect 381154 579978 381774 580046
rect 381154 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 381774 579978
rect 381154 562350 381774 579922
rect 381154 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 381774 562350
rect 381154 562226 381774 562294
rect 381154 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 381774 562226
rect 381154 562102 381774 562170
rect 381154 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 381774 562102
rect 381154 561978 381774 562046
rect 381154 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 381774 561978
rect 381154 544350 381774 561922
rect 381154 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 381774 544350
rect 381154 544226 381774 544294
rect 381154 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 381774 544226
rect 381154 544102 381774 544170
rect 381154 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 381774 544102
rect 381154 543978 381774 544046
rect 381154 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 381774 543978
rect 381154 526350 381774 543922
rect 381154 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 381774 526350
rect 381154 526226 381774 526294
rect 381154 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 381774 526226
rect 381154 526102 381774 526170
rect 381154 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 381774 526102
rect 381154 525978 381774 526046
rect 381154 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 381774 525978
rect 381154 520886 381774 525922
rect 384874 598172 385494 598268
rect 384874 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 385494 598172
rect 384874 598048 385494 598116
rect 384874 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 385494 598048
rect 384874 597924 385494 597992
rect 384874 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 385494 597924
rect 384874 597800 385494 597868
rect 384874 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 385494 597800
rect 384874 586350 385494 597744
rect 384874 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 385494 586350
rect 384874 586226 385494 586294
rect 384874 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 385494 586226
rect 384874 586102 385494 586170
rect 384874 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 385494 586102
rect 384874 585978 385494 586046
rect 384874 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 385494 585978
rect 384874 568350 385494 585922
rect 384874 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 385494 568350
rect 384874 568226 385494 568294
rect 384874 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 385494 568226
rect 384874 568102 385494 568170
rect 384874 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 385494 568102
rect 384874 567978 385494 568046
rect 384874 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 385494 567978
rect 384874 550350 385494 567922
rect 384874 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 385494 550350
rect 384874 550226 385494 550294
rect 384874 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 385494 550226
rect 384874 550102 385494 550170
rect 384874 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 385494 550102
rect 384874 549978 385494 550046
rect 384874 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 385494 549978
rect 384874 532350 385494 549922
rect 384874 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 385494 532350
rect 384874 532226 385494 532294
rect 384874 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 385494 532226
rect 384874 532102 385494 532170
rect 384874 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 385494 532102
rect 384874 531978 385494 532046
rect 384874 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 385494 531978
rect 384874 520886 385494 531922
rect 399154 597212 399774 598268
rect 399154 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 399774 597212
rect 399154 597088 399774 597156
rect 399154 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 399774 597088
rect 399154 596964 399774 597032
rect 399154 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 399774 596964
rect 399154 596840 399774 596908
rect 399154 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 399774 596840
rect 399154 580350 399774 596784
rect 399154 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 399774 580350
rect 399154 580226 399774 580294
rect 399154 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 399774 580226
rect 399154 580102 399774 580170
rect 399154 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 399774 580102
rect 399154 579978 399774 580046
rect 399154 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 399774 579978
rect 399154 562350 399774 579922
rect 399154 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 399774 562350
rect 399154 562226 399774 562294
rect 399154 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 399774 562226
rect 399154 562102 399774 562170
rect 399154 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 399774 562102
rect 399154 561978 399774 562046
rect 399154 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 399774 561978
rect 399154 544350 399774 561922
rect 399154 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 399774 544350
rect 399154 544226 399774 544294
rect 399154 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 399774 544226
rect 399154 544102 399774 544170
rect 399154 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 399774 544102
rect 399154 543978 399774 544046
rect 399154 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 399774 543978
rect 399154 526350 399774 543922
rect 399154 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 399774 526350
rect 399154 526226 399774 526294
rect 399154 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 399774 526226
rect 399154 526102 399774 526170
rect 399154 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 399774 526102
rect 399154 525978 399774 526046
rect 399154 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 399774 525978
rect 399154 520886 399774 525922
rect 402874 598172 403494 598268
rect 402874 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 403494 598172
rect 402874 598048 403494 598116
rect 402874 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 403494 598048
rect 402874 597924 403494 597992
rect 402874 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 403494 597924
rect 402874 597800 403494 597868
rect 402874 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 403494 597800
rect 402874 586350 403494 597744
rect 402874 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 403494 586350
rect 402874 586226 403494 586294
rect 402874 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 403494 586226
rect 402874 586102 403494 586170
rect 402874 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 403494 586102
rect 402874 585978 403494 586046
rect 402874 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 403494 585978
rect 402874 568350 403494 585922
rect 402874 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 403494 568350
rect 402874 568226 403494 568294
rect 402874 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 403494 568226
rect 402874 568102 403494 568170
rect 402874 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 403494 568102
rect 402874 567978 403494 568046
rect 402874 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 403494 567978
rect 402874 550350 403494 567922
rect 402874 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 403494 550350
rect 402874 550226 403494 550294
rect 402874 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 403494 550226
rect 402874 550102 403494 550170
rect 402874 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 403494 550102
rect 402874 549978 403494 550046
rect 402874 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 403494 549978
rect 402874 532350 403494 549922
rect 402874 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 403494 532350
rect 402874 532226 403494 532294
rect 402874 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 403494 532226
rect 402874 532102 403494 532170
rect 402874 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 403494 532102
rect 402874 531978 403494 532046
rect 402874 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 403494 531978
rect 402874 520886 403494 531922
rect 417154 597212 417774 598268
rect 417154 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 417774 597212
rect 417154 597088 417774 597156
rect 417154 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 417774 597088
rect 417154 596964 417774 597032
rect 417154 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 417774 596964
rect 417154 596840 417774 596908
rect 417154 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 417774 596840
rect 417154 580350 417774 596784
rect 417154 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 417774 580350
rect 417154 580226 417774 580294
rect 417154 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 417774 580226
rect 417154 580102 417774 580170
rect 417154 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 417774 580102
rect 417154 579978 417774 580046
rect 417154 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 417774 579978
rect 417154 562350 417774 579922
rect 417154 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 417774 562350
rect 417154 562226 417774 562294
rect 417154 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 417774 562226
rect 417154 562102 417774 562170
rect 417154 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 417774 562102
rect 417154 561978 417774 562046
rect 417154 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 417774 561978
rect 417154 544350 417774 561922
rect 417154 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 417774 544350
rect 417154 544226 417774 544294
rect 417154 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 417774 544226
rect 417154 544102 417774 544170
rect 417154 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 417774 544102
rect 417154 543978 417774 544046
rect 417154 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 417774 543978
rect 417154 526350 417774 543922
rect 417154 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 417774 526350
rect 417154 526226 417774 526294
rect 417154 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 417774 526226
rect 417154 526102 417774 526170
rect 417154 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 417774 526102
rect 417154 525978 417774 526046
rect 417154 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 417774 525978
rect 417154 520886 417774 525922
rect 420874 598172 421494 598268
rect 420874 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 421494 598172
rect 420874 598048 421494 598116
rect 420874 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 421494 598048
rect 420874 597924 421494 597992
rect 420874 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 421494 597924
rect 420874 597800 421494 597868
rect 420874 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 421494 597800
rect 420874 586350 421494 597744
rect 420874 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 421494 586350
rect 420874 586226 421494 586294
rect 420874 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 421494 586226
rect 420874 586102 421494 586170
rect 420874 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 421494 586102
rect 420874 585978 421494 586046
rect 420874 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 421494 585978
rect 420874 568350 421494 585922
rect 420874 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 421494 568350
rect 420874 568226 421494 568294
rect 420874 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 421494 568226
rect 420874 568102 421494 568170
rect 420874 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 421494 568102
rect 420874 567978 421494 568046
rect 420874 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 421494 567978
rect 420874 550350 421494 567922
rect 420874 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 421494 550350
rect 420874 550226 421494 550294
rect 420874 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 421494 550226
rect 420874 550102 421494 550170
rect 420874 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 421494 550102
rect 420874 549978 421494 550046
rect 420874 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 421494 549978
rect 420874 532350 421494 549922
rect 420874 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 421494 532350
rect 420874 532226 421494 532294
rect 420874 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 421494 532226
rect 420874 532102 421494 532170
rect 420874 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 421494 532102
rect 420874 531978 421494 532046
rect 420874 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 421494 531978
rect 420874 520886 421494 531922
rect 435154 597212 435774 598268
rect 435154 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 435774 597212
rect 435154 597088 435774 597156
rect 435154 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 435774 597088
rect 435154 596964 435774 597032
rect 435154 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 435774 596964
rect 435154 596840 435774 596908
rect 435154 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 435774 596840
rect 435154 580350 435774 596784
rect 435154 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 435774 580350
rect 435154 580226 435774 580294
rect 435154 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 435774 580226
rect 435154 580102 435774 580170
rect 435154 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 435774 580102
rect 435154 579978 435774 580046
rect 435154 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 435774 579978
rect 435154 562350 435774 579922
rect 435154 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 435774 562350
rect 435154 562226 435774 562294
rect 435154 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 435774 562226
rect 435154 562102 435774 562170
rect 435154 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 435774 562102
rect 435154 561978 435774 562046
rect 435154 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 435774 561978
rect 435154 544350 435774 561922
rect 435154 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 435774 544350
rect 435154 544226 435774 544294
rect 435154 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 435774 544226
rect 435154 544102 435774 544170
rect 435154 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 435774 544102
rect 435154 543978 435774 544046
rect 435154 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 435774 543978
rect 435154 526350 435774 543922
rect 435154 526294 435250 526350
rect 435306 526294 435374 526350
rect 435430 526294 435498 526350
rect 435554 526294 435622 526350
rect 435678 526294 435774 526350
rect 435154 526226 435774 526294
rect 435154 526170 435250 526226
rect 435306 526170 435374 526226
rect 435430 526170 435498 526226
rect 435554 526170 435622 526226
rect 435678 526170 435774 526226
rect 435154 526102 435774 526170
rect 435154 526046 435250 526102
rect 435306 526046 435374 526102
rect 435430 526046 435498 526102
rect 435554 526046 435622 526102
rect 435678 526046 435774 526102
rect 435154 525978 435774 526046
rect 435154 525922 435250 525978
rect 435306 525922 435374 525978
rect 435430 525922 435498 525978
rect 435554 525922 435622 525978
rect 435678 525922 435774 525978
rect 435154 520886 435774 525922
rect 438874 598172 439494 598268
rect 438874 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 439494 598172
rect 438874 598048 439494 598116
rect 438874 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 439494 598048
rect 438874 597924 439494 597992
rect 438874 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 439494 597924
rect 438874 597800 439494 597868
rect 438874 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 439494 597800
rect 438874 586350 439494 597744
rect 438874 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 439494 586350
rect 438874 586226 439494 586294
rect 438874 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 439494 586226
rect 438874 586102 439494 586170
rect 438874 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 439494 586102
rect 438874 585978 439494 586046
rect 438874 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 439494 585978
rect 438874 568350 439494 585922
rect 438874 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 439494 568350
rect 438874 568226 439494 568294
rect 438874 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 439494 568226
rect 438874 568102 439494 568170
rect 438874 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 439494 568102
rect 438874 567978 439494 568046
rect 438874 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 439494 567978
rect 438874 550350 439494 567922
rect 438874 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 439494 550350
rect 438874 550226 439494 550294
rect 438874 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 439494 550226
rect 438874 550102 439494 550170
rect 438874 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 439494 550102
rect 438874 549978 439494 550046
rect 438874 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 439494 549978
rect 438874 532350 439494 549922
rect 438874 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 439494 532350
rect 438874 532226 439494 532294
rect 438874 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 439494 532226
rect 438874 532102 439494 532170
rect 438874 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 439494 532102
rect 438874 531978 439494 532046
rect 438874 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 439494 531978
rect 438874 520886 439494 531922
rect 453154 597212 453774 598268
rect 453154 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 453774 597212
rect 453154 597088 453774 597156
rect 453154 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 453774 597088
rect 453154 596964 453774 597032
rect 453154 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 453774 596964
rect 453154 596840 453774 596908
rect 453154 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 453774 596840
rect 453154 580350 453774 596784
rect 453154 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 453774 580350
rect 453154 580226 453774 580294
rect 453154 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 453774 580226
rect 453154 580102 453774 580170
rect 453154 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 453774 580102
rect 453154 579978 453774 580046
rect 453154 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 453774 579978
rect 453154 562350 453774 579922
rect 453154 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 453774 562350
rect 453154 562226 453774 562294
rect 453154 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 453774 562226
rect 453154 562102 453774 562170
rect 453154 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 453774 562102
rect 453154 561978 453774 562046
rect 453154 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 453774 561978
rect 453154 544350 453774 561922
rect 453154 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 453774 544350
rect 453154 544226 453774 544294
rect 453154 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 453774 544226
rect 453154 544102 453774 544170
rect 453154 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 453774 544102
rect 453154 543978 453774 544046
rect 453154 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 453774 543978
rect 453154 526350 453774 543922
rect 453154 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 453774 526350
rect 453154 526226 453774 526294
rect 453154 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 453774 526226
rect 453154 526102 453774 526170
rect 453154 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 453774 526102
rect 453154 525978 453774 526046
rect 453154 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 453774 525978
rect 453154 520886 453774 525922
rect 456874 598172 457494 598268
rect 456874 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 457494 598172
rect 456874 598048 457494 598116
rect 456874 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 457494 598048
rect 456874 597924 457494 597992
rect 456874 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 457494 597924
rect 456874 597800 457494 597868
rect 456874 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 457494 597800
rect 456874 586350 457494 597744
rect 456874 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 457494 586350
rect 456874 586226 457494 586294
rect 456874 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 457494 586226
rect 456874 586102 457494 586170
rect 456874 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 457494 586102
rect 456874 585978 457494 586046
rect 456874 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 457494 585978
rect 456874 568350 457494 585922
rect 456874 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 457494 568350
rect 456874 568226 457494 568294
rect 456874 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 457494 568226
rect 456874 568102 457494 568170
rect 456874 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 457494 568102
rect 456874 567978 457494 568046
rect 456874 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 457494 567978
rect 456874 550350 457494 567922
rect 456874 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 457494 550350
rect 456874 550226 457494 550294
rect 456874 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 457494 550226
rect 456874 550102 457494 550170
rect 456874 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 457494 550102
rect 456874 549978 457494 550046
rect 456874 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 457494 549978
rect 456874 532350 457494 549922
rect 456874 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 457494 532350
rect 456874 532226 457494 532294
rect 456874 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 457494 532226
rect 456874 532102 457494 532170
rect 456874 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 457494 532102
rect 456874 531978 457494 532046
rect 456874 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 457494 531978
rect 456874 520886 457494 531922
rect 471154 597212 471774 598268
rect 471154 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 471774 597212
rect 471154 597088 471774 597156
rect 471154 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 471774 597088
rect 471154 596964 471774 597032
rect 471154 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 471774 596964
rect 471154 596840 471774 596908
rect 471154 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 471774 596840
rect 471154 580350 471774 596784
rect 471154 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 471774 580350
rect 471154 580226 471774 580294
rect 471154 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 471774 580226
rect 471154 580102 471774 580170
rect 471154 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 471774 580102
rect 471154 579978 471774 580046
rect 471154 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 471774 579978
rect 471154 562350 471774 579922
rect 471154 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 471774 562350
rect 471154 562226 471774 562294
rect 471154 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 471774 562226
rect 471154 562102 471774 562170
rect 471154 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 471774 562102
rect 471154 561978 471774 562046
rect 471154 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 471774 561978
rect 471154 544350 471774 561922
rect 471154 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 471774 544350
rect 471154 544226 471774 544294
rect 471154 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 471774 544226
rect 471154 544102 471774 544170
rect 471154 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 471774 544102
rect 471154 543978 471774 544046
rect 471154 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 471774 543978
rect 471154 526350 471774 543922
rect 471154 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 471774 526350
rect 471154 526226 471774 526294
rect 471154 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 471774 526226
rect 471154 526102 471774 526170
rect 471154 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 471774 526102
rect 471154 525978 471774 526046
rect 471154 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 471774 525978
rect 471154 520886 471774 525922
rect 474874 598172 475494 598268
rect 474874 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 475494 598172
rect 474874 598048 475494 598116
rect 474874 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 475494 598048
rect 474874 597924 475494 597992
rect 474874 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 475494 597924
rect 474874 597800 475494 597868
rect 474874 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 475494 597800
rect 474874 586350 475494 597744
rect 474874 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 475494 586350
rect 474874 586226 475494 586294
rect 474874 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 475494 586226
rect 474874 586102 475494 586170
rect 474874 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 475494 586102
rect 474874 585978 475494 586046
rect 474874 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 475494 585978
rect 474874 568350 475494 585922
rect 474874 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 475494 568350
rect 474874 568226 475494 568294
rect 474874 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 475494 568226
rect 474874 568102 475494 568170
rect 474874 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 475494 568102
rect 474874 567978 475494 568046
rect 474874 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 475494 567978
rect 474874 550350 475494 567922
rect 474874 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 475494 550350
rect 474874 550226 475494 550294
rect 474874 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 475494 550226
rect 474874 550102 475494 550170
rect 474874 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 475494 550102
rect 474874 549978 475494 550046
rect 474874 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 475494 549978
rect 474874 532350 475494 549922
rect 474874 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 475494 532350
rect 474874 532226 475494 532294
rect 474874 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 475494 532226
rect 474874 532102 475494 532170
rect 474874 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 475494 532102
rect 474874 531978 475494 532046
rect 474874 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 475494 531978
rect 474874 520886 475494 531922
rect 489154 597212 489774 598268
rect 489154 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 489774 597212
rect 489154 597088 489774 597156
rect 489154 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 489774 597088
rect 489154 596964 489774 597032
rect 489154 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 489774 596964
rect 489154 596840 489774 596908
rect 489154 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 489774 596840
rect 489154 580350 489774 596784
rect 489154 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 489774 580350
rect 489154 580226 489774 580294
rect 489154 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 489774 580226
rect 489154 580102 489774 580170
rect 489154 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 489774 580102
rect 489154 579978 489774 580046
rect 489154 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 489774 579978
rect 489154 562350 489774 579922
rect 489154 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 489774 562350
rect 489154 562226 489774 562294
rect 489154 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 489774 562226
rect 489154 562102 489774 562170
rect 489154 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 489774 562102
rect 489154 561978 489774 562046
rect 489154 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 489774 561978
rect 489154 544350 489774 561922
rect 489154 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 489774 544350
rect 489154 544226 489774 544294
rect 489154 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 489774 544226
rect 489154 544102 489774 544170
rect 489154 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 489774 544102
rect 489154 543978 489774 544046
rect 489154 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 489774 543978
rect 489154 526350 489774 543922
rect 489154 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 489774 526350
rect 489154 526226 489774 526294
rect 489154 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 489774 526226
rect 489154 526102 489774 526170
rect 489154 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 489774 526102
rect 489154 525978 489774 526046
rect 489154 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 489774 525978
rect 489154 520886 489774 525922
rect 492874 598172 493494 598268
rect 492874 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 493494 598172
rect 492874 598048 493494 598116
rect 492874 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 493494 598048
rect 492874 597924 493494 597992
rect 492874 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 493494 597924
rect 492874 597800 493494 597868
rect 492874 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 493494 597800
rect 492874 586350 493494 597744
rect 492874 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 493494 586350
rect 492874 586226 493494 586294
rect 492874 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 493494 586226
rect 492874 586102 493494 586170
rect 492874 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 493494 586102
rect 492874 585978 493494 586046
rect 492874 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 493494 585978
rect 492874 568350 493494 585922
rect 492874 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 493494 568350
rect 492874 568226 493494 568294
rect 492874 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 493494 568226
rect 492874 568102 493494 568170
rect 492874 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 493494 568102
rect 492874 567978 493494 568046
rect 492874 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 493494 567978
rect 492874 550350 493494 567922
rect 492874 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 493494 550350
rect 492874 550226 493494 550294
rect 492874 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 493494 550226
rect 492874 550102 493494 550170
rect 492874 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 493494 550102
rect 492874 549978 493494 550046
rect 492874 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 493494 549978
rect 492874 532350 493494 549922
rect 492874 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 493494 532350
rect 492874 532226 493494 532294
rect 492874 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 493494 532226
rect 492874 532102 493494 532170
rect 492874 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 493494 532102
rect 492874 531978 493494 532046
rect 492874 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 493494 531978
rect 492874 520886 493494 531922
rect 507154 597212 507774 598268
rect 507154 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 507774 597212
rect 507154 597088 507774 597156
rect 507154 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 507774 597088
rect 507154 596964 507774 597032
rect 507154 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 507774 596964
rect 507154 596840 507774 596908
rect 507154 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 507774 596840
rect 507154 580350 507774 596784
rect 507154 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 507774 580350
rect 507154 580226 507774 580294
rect 507154 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 507774 580226
rect 507154 580102 507774 580170
rect 507154 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 507774 580102
rect 507154 579978 507774 580046
rect 507154 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 507774 579978
rect 507154 562350 507774 579922
rect 507154 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 507774 562350
rect 507154 562226 507774 562294
rect 507154 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 507774 562226
rect 507154 562102 507774 562170
rect 507154 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 507774 562102
rect 507154 561978 507774 562046
rect 507154 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 507774 561978
rect 507154 544350 507774 561922
rect 507154 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 507774 544350
rect 507154 544226 507774 544294
rect 507154 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 507774 544226
rect 507154 544102 507774 544170
rect 507154 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 507774 544102
rect 507154 543978 507774 544046
rect 507154 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 507774 543978
rect 507154 526350 507774 543922
rect 507154 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 507774 526350
rect 507154 526226 507774 526294
rect 507154 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 507774 526226
rect 507154 526102 507774 526170
rect 507154 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 507774 526102
rect 507154 525978 507774 526046
rect 507154 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 507774 525978
rect 507154 520886 507774 525922
rect 510874 598172 511494 598268
rect 510874 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 511494 598172
rect 510874 598048 511494 598116
rect 510874 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 511494 598048
rect 510874 597924 511494 597992
rect 510874 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 511494 597924
rect 510874 597800 511494 597868
rect 510874 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 511494 597800
rect 510874 586350 511494 597744
rect 510874 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 511494 586350
rect 510874 586226 511494 586294
rect 510874 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 511494 586226
rect 510874 586102 511494 586170
rect 510874 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 511494 586102
rect 510874 585978 511494 586046
rect 510874 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 511494 585978
rect 510874 568350 511494 585922
rect 510874 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 511494 568350
rect 510874 568226 511494 568294
rect 510874 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 511494 568226
rect 510874 568102 511494 568170
rect 510874 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 511494 568102
rect 510874 567978 511494 568046
rect 510874 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 511494 567978
rect 510874 550350 511494 567922
rect 510874 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 511494 550350
rect 510874 550226 511494 550294
rect 510874 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 511494 550226
rect 510874 550102 511494 550170
rect 510874 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 511494 550102
rect 510874 549978 511494 550046
rect 510874 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 511494 549978
rect 510874 532350 511494 549922
rect 510874 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 511494 532350
rect 510874 532226 511494 532294
rect 510874 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 511494 532226
rect 510874 532102 511494 532170
rect 510874 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 511494 532102
rect 510874 531978 511494 532046
rect 510874 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 511494 531978
rect 510874 520886 511494 531922
rect 525154 597212 525774 598268
rect 525154 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 525774 597212
rect 525154 597088 525774 597156
rect 525154 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 525774 597088
rect 525154 596964 525774 597032
rect 525154 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 525774 596964
rect 525154 596840 525774 596908
rect 525154 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 525774 596840
rect 525154 580350 525774 596784
rect 525154 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 525774 580350
rect 525154 580226 525774 580294
rect 525154 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 525774 580226
rect 525154 580102 525774 580170
rect 525154 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 525774 580102
rect 525154 579978 525774 580046
rect 525154 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 525774 579978
rect 525154 562350 525774 579922
rect 525154 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 525774 562350
rect 525154 562226 525774 562294
rect 525154 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 525774 562226
rect 525154 562102 525774 562170
rect 525154 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 525774 562102
rect 525154 561978 525774 562046
rect 525154 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 525774 561978
rect 525154 544350 525774 561922
rect 525154 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 525774 544350
rect 525154 544226 525774 544294
rect 525154 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 525774 544226
rect 525154 544102 525774 544170
rect 525154 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 525774 544102
rect 525154 543978 525774 544046
rect 525154 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 525774 543978
rect 525154 526350 525774 543922
rect 525154 526294 525250 526350
rect 525306 526294 525374 526350
rect 525430 526294 525498 526350
rect 525554 526294 525622 526350
rect 525678 526294 525774 526350
rect 525154 526226 525774 526294
rect 525154 526170 525250 526226
rect 525306 526170 525374 526226
rect 525430 526170 525498 526226
rect 525554 526170 525622 526226
rect 525678 526170 525774 526226
rect 525154 526102 525774 526170
rect 525154 526046 525250 526102
rect 525306 526046 525374 526102
rect 525430 526046 525498 526102
rect 525554 526046 525622 526102
rect 525678 526046 525774 526102
rect 525154 525978 525774 526046
rect 525154 525922 525250 525978
rect 525306 525922 525374 525978
rect 525430 525922 525498 525978
rect 525554 525922 525622 525978
rect 525678 525922 525774 525978
rect 6874 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 7494 514350
rect 6874 514226 7494 514294
rect 6874 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 7494 514226
rect 6874 514102 7494 514170
rect 6874 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 7494 514102
rect 6874 513978 7494 514046
rect 6874 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 7494 513978
rect 6874 496350 7494 513922
rect 39808 514350 40128 514384
rect 39808 514294 39878 514350
rect 39934 514294 40002 514350
rect 40058 514294 40128 514350
rect 39808 514226 40128 514294
rect 39808 514170 39878 514226
rect 39934 514170 40002 514226
rect 40058 514170 40128 514226
rect 39808 514102 40128 514170
rect 39808 514046 39878 514102
rect 39934 514046 40002 514102
rect 40058 514046 40128 514102
rect 39808 513978 40128 514046
rect 39808 513922 39878 513978
rect 39934 513922 40002 513978
rect 40058 513922 40128 513978
rect 39808 513888 40128 513922
rect 70528 514350 70848 514384
rect 70528 514294 70598 514350
rect 70654 514294 70722 514350
rect 70778 514294 70848 514350
rect 70528 514226 70848 514294
rect 70528 514170 70598 514226
rect 70654 514170 70722 514226
rect 70778 514170 70848 514226
rect 70528 514102 70848 514170
rect 70528 514046 70598 514102
rect 70654 514046 70722 514102
rect 70778 514046 70848 514102
rect 70528 513978 70848 514046
rect 70528 513922 70598 513978
rect 70654 513922 70722 513978
rect 70778 513922 70848 513978
rect 70528 513888 70848 513922
rect 101248 514350 101568 514384
rect 101248 514294 101318 514350
rect 101374 514294 101442 514350
rect 101498 514294 101568 514350
rect 101248 514226 101568 514294
rect 101248 514170 101318 514226
rect 101374 514170 101442 514226
rect 101498 514170 101568 514226
rect 101248 514102 101568 514170
rect 101248 514046 101318 514102
rect 101374 514046 101442 514102
rect 101498 514046 101568 514102
rect 101248 513978 101568 514046
rect 101248 513922 101318 513978
rect 101374 513922 101442 513978
rect 101498 513922 101568 513978
rect 101248 513888 101568 513922
rect 131968 514350 132288 514384
rect 131968 514294 132038 514350
rect 132094 514294 132162 514350
rect 132218 514294 132288 514350
rect 131968 514226 132288 514294
rect 131968 514170 132038 514226
rect 132094 514170 132162 514226
rect 132218 514170 132288 514226
rect 131968 514102 132288 514170
rect 131968 514046 132038 514102
rect 132094 514046 132162 514102
rect 132218 514046 132288 514102
rect 131968 513978 132288 514046
rect 131968 513922 132038 513978
rect 132094 513922 132162 513978
rect 132218 513922 132288 513978
rect 131968 513888 132288 513922
rect 162688 514350 163008 514384
rect 162688 514294 162758 514350
rect 162814 514294 162882 514350
rect 162938 514294 163008 514350
rect 162688 514226 163008 514294
rect 162688 514170 162758 514226
rect 162814 514170 162882 514226
rect 162938 514170 163008 514226
rect 162688 514102 163008 514170
rect 162688 514046 162758 514102
rect 162814 514046 162882 514102
rect 162938 514046 163008 514102
rect 162688 513978 163008 514046
rect 162688 513922 162758 513978
rect 162814 513922 162882 513978
rect 162938 513922 163008 513978
rect 162688 513888 163008 513922
rect 193408 514350 193728 514384
rect 193408 514294 193478 514350
rect 193534 514294 193602 514350
rect 193658 514294 193728 514350
rect 193408 514226 193728 514294
rect 193408 514170 193478 514226
rect 193534 514170 193602 514226
rect 193658 514170 193728 514226
rect 193408 514102 193728 514170
rect 193408 514046 193478 514102
rect 193534 514046 193602 514102
rect 193658 514046 193728 514102
rect 193408 513978 193728 514046
rect 193408 513922 193478 513978
rect 193534 513922 193602 513978
rect 193658 513922 193728 513978
rect 193408 513888 193728 513922
rect 224128 514350 224448 514384
rect 224128 514294 224198 514350
rect 224254 514294 224322 514350
rect 224378 514294 224448 514350
rect 224128 514226 224448 514294
rect 224128 514170 224198 514226
rect 224254 514170 224322 514226
rect 224378 514170 224448 514226
rect 224128 514102 224448 514170
rect 224128 514046 224198 514102
rect 224254 514046 224322 514102
rect 224378 514046 224448 514102
rect 224128 513978 224448 514046
rect 224128 513922 224198 513978
rect 224254 513922 224322 513978
rect 224378 513922 224448 513978
rect 224128 513888 224448 513922
rect 254848 514350 255168 514384
rect 254848 514294 254918 514350
rect 254974 514294 255042 514350
rect 255098 514294 255168 514350
rect 254848 514226 255168 514294
rect 254848 514170 254918 514226
rect 254974 514170 255042 514226
rect 255098 514170 255168 514226
rect 254848 514102 255168 514170
rect 254848 514046 254918 514102
rect 254974 514046 255042 514102
rect 255098 514046 255168 514102
rect 254848 513978 255168 514046
rect 254848 513922 254918 513978
rect 254974 513922 255042 513978
rect 255098 513922 255168 513978
rect 254848 513888 255168 513922
rect 285568 514350 285888 514384
rect 285568 514294 285638 514350
rect 285694 514294 285762 514350
rect 285818 514294 285888 514350
rect 285568 514226 285888 514294
rect 285568 514170 285638 514226
rect 285694 514170 285762 514226
rect 285818 514170 285888 514226
rect 285568 514102 285888 514170
rect 285568 514046 285638 514102
rect 285694 514046 285762 514102
rect 285818 514046 285888 514102
rect 285568 513978 285888 514046
rect 285568 513922 285638 513978
rect 285694 513922 285762 513978
rect 285818 513922 285888 513978
rect 285568 513888 285888 513922
rect 316288 514350 316608 514384
rect 316288 514294 316358 514350
rect 316414 514294 316482 514350
rect 316538 514294 316608 514350
rect 316288 514226 316608 514294
rect 316288 514170 316358 514226
rect 316414 514170 316482 514226
rect 316538 514170 316608 514226
rect 316288 514102 316608 514170
rect 316288 514046 316358 514102
rect 316414 514046 316482 514102
rect 316538 514046 316608 514102
rect 316288 513978 316608 514046
rect 316288 513922 316358 513978
rect 316414 513922 316482 513978
rect 316538 513922 316608 513978
rect 316288 513888 316608 513922
rect 347008 514350 347328 514384
rect 347008 514294 347078 514350
rect 347134 514294 347202 514350
rect 347258 514294 347328 514350
rect 347008 514226 347328 514294
rect 347008 514170 347078 514226
rect 347134 514170 347202 514226
rect 347258 514170 347328 514226
rect 347008 514102 347328 514170
rect 347008 514046 347078 514102
rect 347134 514046 347202 514102
rect 347258 514046 347328 514102
rect 347008 513978 347328 514046
rect 347008 513922 347078 513978
rect 347134 513922 347202 513978
rect 347258 513922 347328 513978
rect 347008 513888 347328 513922
rect 377728 514350 378048 514384
rect 377728 514294 377798 514350
rect 377854 514294 377922 514350
rect 377978 514294 378048 514350
rect 377728 514226 378048 514294
rect 377728 514170 377798 514226
rect 377854 514170 377922 514226
rect 377978 514170 378048 514226
rect 377728 514102 378048 514170
rect 377728 514046 377798 514102
rect 377854 514046 377922 514102
rect 377978 514046 378048 514102
rect 377728 513978 378048 514046
rect 377728 513922 377798 513978
rect 377854 513922 377922 513978
rect 377978 513922 378048 513978
rect 377728 513888 378048 513922
rect 408448 514350 408768 514384
rect 408448 514294 408518 514350
rect 408574 514294 408642 514350
rect 408698 514294 408768 514350
rect 408448 514226 408768 514294
rect 408448 514170 408518 514226
rect 408574 514170 408642 514226
rect 408698 514170 408768 514226
rect 408448 514102 408768 514170
rect 408448 514046 408518 514102
rect 408574 514046 408642 514102
rect 408698 514046 408768 514102
rect 408448 513978 408768 514046
rect 408448 513922 408518 513978
rect 408574 513922 408642 513978
rect 408698 513922 408768 513978
rect 408448 513888 408768 513922
rect 439168 514350 439488 514384
rect 439168 514294 439238 514350
rect 439294 514294 439362 514350
rect 439418 514294 439488 514350
rect 439168 514226 439488 514294
rect 439168 514170 439238 514226
rect 439294 514170 439362 514226
rect 439418 514170 439488 514226
rect 439168 514102 439488 514170
rect 439168 514046 439238 514102
rect 439294 514046 439362 514102
rect 439418 514046 439488 514102
rect 439168 513978 439488 514046
rect 439168 513922 439238 513978
rect 439294 513922 439362 513978
rect 439418 513922 439488 513978
rect 439168 513888 439488 513922
rect 469888 514350 470208 514384
rect 469888 514294 469958 514350
rect 470014 514294 470082 514350
rect 470138 514294 470208 514350
rect 469888 514226 470208 514294
rect 469888 514170 469958 514226
rect 470014 514170 470082 514226
rect 470138 514170 470208 514226
rect 469888 514102 470208 514170
rect 469888 514046 469958 514102
rect 470014 514046 470082 514102
rect 470138 514046 470208 514102
rect 469888 513978 470208 514046
rect 469888 513922 469958 513978
rect 470014 513922 470082 513978
rect 470138 513922 470208 513978
rect 469888 513888 470208 513922
rect 500608 514350 500928 514384
rect 500608 514294 500678 514350
rect 500734 514294 500802 514350
rect 500858 514294 500928 514350
rect 500608 514226 500928 514294
rect 500608 514170 500678 514226
rect 500734 514170 500802 514226
rect 500858 514170 500928 514226
rect 500608 514102 500928 514170
rect 500608 514046 500678 514102
rect 500734 514046 500802 514102
rect 500858 514046 500928 514102
rect 500608 513978 500928 514046
rect 500608 513922 500678 513978
rect 500734 513922 500802 513978
rect 500858 513922 500928 513978
rect 500608 513888 500928 513922
rect 24448 508350 24768 508384
rect 24448 508294 24518 508350
rect 24574 508294 24642 508350
rect 24698 508294 24768 508350
rect 24448 508226 24768 508294
rect 24448 508170 24518 508226
rect 24574 508170 24642 508226
rect 24698 508170 24768 508226
rect 24448 508102 24768 508170
rect 24448 508046 24518 508102
rect 24574 508046 24642 508102
rect 24698 508046 24768 508102
rect 24448 507978 24768 508046
rect 24448 507922 24518 507978
rect 24574 507922 24642 507978
rect 24698 507922 24768 507978
rect 24448 507888 24768 507922
rect 55168 508350 55488 508384
rect 55168 508294 55238 508350
rect 55294 508294 55362 508350
rect 55418 508294 55488 508350
rect 55168 508226 55488 508294
rect 55168 508170 55238 508226
rect 55294 508170 55362 508226
rect 55418 508170 55488 508226
rect 55168 508102 55488 508170
rect 55168 508046 55238 508102
rect 55294 508046 55362 508102
rect 55418 508046 55488 508102
rect 55168 507978 55488 508046
rect 55168 507922 55238 507978
rect 55294 507922 55362 507978
rect 55418 507922 55488 507978
rect 55168 507888 55488 507922
rect 85888 508350 86208 508384
rect 85888 508294 85958 508350
rect 86014 508294 86082 508350
rect 86138 508294 86208 508350
rect 85888 508226 86208 508294
rect 85888 508170 85958 508226
rect 86014 508170 86082 508226
rect 86138 508170 86208 508226
rect 85888 508102 86208 508170
rect 85888 508046 85958 508102
rect 86014 508046 86082 508102
rect 86138 508046 86208 508102
rect 85888 507978 86208 508046
rect 85888 507922 85958 507978
rect 86014 507922 86082 507978
rect 86138 507922 86208 507978
rect 85888 507888 86208 507922
rect 116608 508350 116928 508384
rect 116608 508294 116678 508350
rect 116734 508294 116802 508350
rect 116858 508294 116928 508350
rect 116608 508226 116928 508294
rect 116608 508170 116678 508226
rect 116734 508170 116802 508226
rect 116858 508170 116928 508226
rect 116608 508102 116928 508170
rect 116608 508046 116678 508102
rect 116734 508046 116802 508102
rect 116858 508046 116928 508102
rect 116608 507978 116928 508046
rect 116608 507922 116678 507978
rect 116734 507922 116802 507978
rect 116858 507922 116928 507978
rect 116608 507888 116928 507922
rect 147328 508350 147648 508384
rect 147328 508294 147398 508350
rect 147454 508294 147522 508350
rect 147578 508294 147648 508350
rect 147328 508226 147648 508294
rect 147328 508170 147398 508226
rect 147454 508170 147522 508226
rect 147578 508170 147648 508226
rect 147328 508102 147648 508170
rect 147328 508046 147398 508102
rect 147454 508046 147522 508102
rect 147578 508046 147648 508102
rect 147328 507978 147648 508046
rect 147328 507922 147398 507978
rect 147454 507922 147522 507978
rect 147578 507922 147648 507978
rect 147328 507888 147648 507922
rect 178048 508350 178368 508384
rect 178048 508294 178118 508350
rect 178174 508294 178242 508350
rect 178298 508294 178368 508350
rect 178048 508226 178368 508294
rect 178048 508170 178118 508226
rect 178174 508170 178242 508226
rect 178298 508170 178368 508226
rect 178048 508102 178368 508170
rect 178048 508046 178118 508102
rect 178174 508046 178242 508102
rect 178298 508046 178368 508102
rect 178048 507978 178368 508046
rect 178048 507922 178118 507978
rect 178174 507922 178242 507978
rect 178298 507922 178368 507978
rect 178048 507888 178368 507922
rect 208768 508350 209088 508384
rect 208768 508294 208838 508350
rect 208894 508294 208962 508350
rect 209018 508294 209088 508350
rect 208768 508226 209088 508294
rect 208768 508170 208838 508226
rect 208894 508170 208962 508226
rect 209018 508170 209088 508226
rect 208768 508102 209088 508170
rect 208768 508046 208838 508102
rect 208894 508046 208962 508102
rect 209018 508046 209088 508102
rect 208768 507978 209088 508046
rect 208768 507922 208838 507978
rect 208894 507922 208962 507978
rect 209018 507922 209088 507978
rect 208768 507888 209088 507922
rect 239488 508350 239808 508384
rect 239488 508294 239558 508350
rect 239614 508294 239682 508350
rect 239738 508294 239808 508350
rect 239488 508226 239808 508294
rect 239488 508170 239558 508226
rect 239614 508170 239682 508226
rect 239738 508170 239808 508226
rect 239488 508102 239808 508170
rect 239488 508046 239558 508102
rect 239614 508046 239682 508102
rect 239738 508046 239808 508102
rect 239488 507978 239808 508046
rect 239488 507922 239558 507978
rect 239614 507922 239682 507978
rect 239738 507922 239808 507978
rect 239488 507888 239808 507922
rect 270208 508350 270528 508384
rect 270208 508294 270278 508350
rect 270334 508294 270402 508350
rect 270458 508294 270528 508350
rect 270208 508226 270528 508294
rect 270208 508170 270278 508226
rect 270334 508170 270402 508226
rect 270458 508170 270528 508226
rect 270208 508102 270528 508170
rect 270208 508046 270278 508102
rect 270334 508046 270402 508102
rect 270458 508046 270528 508102
rect 270208 507978 270528 508046
rect 270208 507922 270278 507978
rect 270334 507922 270402 507978
rect 270458 507922 270528 507978
rect 270208 507888 270528 507922
rect 300928 508350 301248 508384
rect 300928 508294 300998 508350
rect 301054 508294 301122 508350
rect 301178 508294 301248 508350
rect 300928 508226 301248 508294
rect 300928 508170 300998 508226
rect 301054 508170 301122 508226
rect 301178 508170 301248 508226
rect 300928 508102 301248 508170
rect 300928 508046 300998 508102
rect 301054 508046 301122 508102
rect 301178 508046 301248 508102
rect 300928 507978 301248 508046
rect 300928 507922 300998 507978
rect 301054 507922 301122 507978
rect 301178 507922 301248 507978
rect 300928 507888 301248 507922
rect 331648 508350 331968 508384
rect 331648 508294 331718 508350
rect 331774 508294 331842 508350
rect 331898 508294 331968 508350
rect 331648 508226 331968 508294
rect 331648 508170 331718 508226
rect 331774 508170 331842 508226
rect 331898 508170 331968 508226
rect 331648 508102 331968 508170
rect 331648 508046 331718 508102
rect 331774 508046 331842 508102
rect 331898 508046 331968 508102
rect 331648 507978 331968 508046
rect 331648 507922 331718 507978
rect 331774 507922 331842 507978
rect 331898 507922 331968 507978
rect 331648 507888 331968 507922
rect 362368 508350 362688 508384
rect 362368 508294 362438 508350
rect 362494 508294 362562 508350
rect 362618 508294 362688 508350
rect 362368 508226 362688 508294
rect 362368 508170 362438 508226
rect 362494 508170 362562 508226
rect 362618 508170 362688 508226
rect 362368 508102 362688 508170
rect 362368 508046 362438 508102
rect 362494 508046 362562 508102
rect 362618 508046 362688 508102
rect 362368 507978 362688 508046
rect 362368 507922 362438 507978
rect 362494 507922 362562 507978
rect 362618 507922 362688 507978
rect 362368 507888 362688 507922
rect 393088 508350 393408 508384
rect 393088 508294 393158 508350
rect 393214 508294 393282 508350
rect 393338 508294 393408 508350
rect 393088 508226 393408 508294
rect 393088 508170 393158 508226
rect 393214 508170 393282 508226
rect 393338 508170 393408 508226
rect 393088 508102 393408 508170
rect 393088 508046 393158 508102
rect 393214 508046 393282 508102
rect 393338 508046 393408 508102
rect 393088 507978 393408 508046
rect 393088 507922 393158 507978
rect 393214 507922 393282 507978
rect 393338 507922 393408 507978
rect 393088 507888 393408 507922
rect 423808 508350 424128 508384
rect 423808 508294 423878 508350
rect 423934 508294 424002 508350
rect 424058 508294 424128 508350
rect 423808 508226 424128 508294
rect 423808 508170 423878 508226
rect 423934 508170 424002 508226
rect 424058 508170 424128 508226
rect 423808 508102 424128 508170
rect 423808 508046 423878 508102
rect 423934 508046 424002 508102
rect 424058 508046 424128 508102
rect 423808 507978 424128 508046
rect 423808 507922 423878 507978
rect 423934 507922 424002 507978
rect 424058 507922 424128 507978
rect 423808 507888 424128 507922
rect 454528 508350 454848 508384
rect 454528 508294 454598 508350
rect 454654 508294 454722 508350
rect 454778 508294 454848 508350
rect 454528 508226 454848 508294
rect 454528 508170 454598 508226
rect 454654 508170 454722 508226
rect 454778 508170 454848 508226
rect 454528 508102 454848 508170
rect 454528 508046 454598 508102
rect 454654 508046 454722 508102
rect 454778 508046 454848 508102
rect 454528 507978 454848 508046
rect 454528 507922 454598 507978
rect 454654 507922 454722 507978
rect 454778 507922 454848 507978
rect 454528 507888 454848 507922
rect 485248 508350 485568 508384
rect 485248 508294 485318 508350
rect 485374 508294 485442 508350
rect 485498 508294 485568 508350
rect 485248 508226 485568 508294
rect 485248 508170 485318 508226
rect 485374 508170 485442 508226
rect 485498 508170 485568 508226
rect 485248 508102 485568 508170
rect 485248 508046 485318 508102
rect 485374 508046 485442 508102
rect 485498 508046 485568 508102
rect 485248 507978 485568 508046
rect 485248 507922 485318 507978
rect 485374 507922 485442 507978
rect 485498 507922 485568 507978
rect 485248 507888 485568 507922
rect 515968 508350 516288 508384
rect 515968 508294 516038 508350
rect 516094 508294 516162 508350
rect 516218 508294 516288 508350
rect 515968 508226 516288 508294
rect 515968 508170 516038 508226
rect 516094 508170 516162 508226
rect 516218 508170 516288 508226
rect 515968 508102 516288 508170
rect 515968 508046 516038 508102
rect 516094 508046 516162 508102
rect 516218 508046 516288 508102
rect 515968 507978 516288 508046
rect 515968 507922 516038 507978
rect 516094 507922 516162 507978
rect 516218 507922 516288 507978
rect 515968 507888 516288 507922
rect 525154 508350 525774 525922
rect 525154 508294 525250 508350
rect 525306 508294 525374 508350
rect 525430 508294 525498 508350
rect 525554 508294 525622 508350
rect 525678 508294 525774 508350
rect 525154 508226 525774 508294
rect 525154 508170 525250 508226
rect 525306 508170 525374 508226
rect 525430 508170 525498 508226
rect 525554 508170 525622 508226
rect 525678 508170 525774 508226
rect 525154 508102 525774 508170
rect 525154 508046 525250 508102
rect 525306 508046 525374 508102
rect 525430 508046 525498 508102
rect 525554 508046 525622 508102
rect 525678 508046 525774 508102
rect 525154 507978 525774 508046
rect 525154 507922 525250 507978
rect 525306 507922 525374 507978
rect 525430 507922 525498 507978
rect 525554 507922 525622 507978
rect 525678 507922 525774 507978
rect 6874 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 7494 496350
rect 6874 496226 7494 496294
rect 6874 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 7494 496226
rect 6874 496102 7494 496170
rect 6874 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 7494 496102
rect 6874 495978 7494 496046
rect 6874 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 7494 495978
rect 6874 478350 7494 495922
rect 39808 496350 40128 496384
rect 39808 496294 39878 496350
rect 39934 496294 40002 496350
rect 40058 496294 40128 496350
rect 39808 496226 40128 496294
rect 39808 496170 39878 496226
rect 39934 496170 40002 496226
rect 40058 496170 40128 496226
rect 39808 496102 40128 496170
rect 39808 496046 39878 496102
rect 39934 496046 40002 496102
rect 40058 496046 40128 496102
rect 39808 495978 40128 496046
rect 39808 495922 39878 495978
rect 39934 495922 40002 495978
rect 40058 495922 40128 495978
rect 39808 495888 40128 495922
rect 70528 496350 70848 496384
rect 70528 496294 70598 496350
rect 70654 496294 70722 496350
rect 70778 496294 70848 496350
rect 70528 496226 70848 496294
rect 70528 496170 70598 496226
rect 70654 496170 70722 496226
rect 70778 496170 70848 496226
rect 70528 496102 70848 496170
rect 70528 496046 70598 496102
rect 70654 496046 70722 496102
rect 70778 496046 70848 496102
rect 70528 495978 70848 496046
rect 70528 495922 70598 495978
rect 70654 495922 70722 495978
rect 70778 495922 70848 495978
rect 70528 495888 70848 495922
rect 101248 496350 101568 496384
rect 101248 496294 101318 496350
rect 101374 496294 101442 496350
rect 101498 496294 101568 496350
rect 101248 496226 101568 496294
rect 101248 496170 101318 496226
rect 101374 496170 101442 496226
rect 101498 496170 101568 496226
rect 101248 496102 101568 496170
rect 101248 496046 101318 496102
rect 101374 496046 101442 496102
rect 101498 496046 101568 496102
rect 101248 495978 101568 496046
rect 101248 495922 101318 495978
rect 101374 495922 101442 495978
rect 101498 495922 101568 495978
rect 101248 495888 101568 495922
rect 131968 496350 132288 496384
rect 131968 496294 132038 496350
rect 132094 496294 132162 496350
rect 132218 496294 132288 496350
rect 131968 496226 132288 496294
rect 131968 496170 132038 496226
rect 132094 496170 132162 496226
rect 132218 496170 132288 496226
rect 131968 496102 132288 496170
rect 131968 496046 132038 496102
rect 132094 496046 132162 496102
rect 132218 496046 132288 496102
rect 131968 495978 132288 496046
rect 131968 495922 132038 495978
rect 132094 495922 132162 495978
rect 132218 495922 132288 495978
rect 131968 495888 132288 495922
rect 162688 496350 163008 496384
rect 162688 496294 162758 496350
rect 162814 496294 162882 496350
rect 162938 496294 163008 496350
rect 162688 496226 163008 496294
rect 162688 496170 162758 496226
rect 162814 496170 162882 496226
rect 162938 496170 163008 496226
rect 162688 496102 163008 496170
rect 162688 496046 162758 496102
rect 162814 496046 162882 496102
rect 162938 496046 163008 496102
rect 162688 495978 163008 496046
rect 162688 495922 162758 495978
rect 162814 495922 162882 495978
rect 162938 495922 163008 495978
rect 162688 495888 163008 495922
rect 193408 496350 193728 496384
rect 193408 496294 193478 496350
rect 193534 496294 193602 496350
rect 193658 496294 193728 496350
rect 193408 496226 193728 496294
rect 193408 496170 193478 496226
rect 193534 496170 193602 496226
rect 193658 496170 193728 496226
rect 193408 496102 193728 496170
rect 193408 496046 193478 496102
rect 193534 496046 193602 496102
rect 193658 496046 193728 496102
rect 193408 495978 193728 496046
rect 193408 495922 193478 495978
rect 193534 495922 193602 495978
rect 193658 495922 193728 495978
rect 193408 495888 193728 495922
rect 224128 496350 224448 496384
rect 224128 496294 224198 496350
rect 224254 496294 224322 496350
rect 224378 496294 224448 496350
rect 224128 496226 224448 496294
rect 224128 496170 224198 496226
rect 224254 496170 224322 496226
rect 224378 496170 224448 496226
rect 224128 496102 224448 496170
rect 224128 496046 224198 496102
rect 224254 496046 224322 496102
rect 224378 496046 224448 496102
rect 224128 495978 224448 496046
rect 224128 495922 224198 495978
rect 224254 495922 224322 495978
rect 224378 495922 224448 495978
rect 224128 495888 224448 495922
rect 254848 496350 255168 496384
rect 254848 496294 254918 496350
rect 254974 496294 255042 496350
rect 255098 496294 255168 496350
rect 254848 496226 255168 496294
rect 254848 496170 254918 496226
rect 254974 496170 255042 496226
rect 255098 496170 255168 496226
rect 254848 496102 255168 496170
rect 254848 496046 254918 496102
rect 254974 496046 255042 496102
rect 255098 496046 255168 496102
rect 254848 495978 255168 496046
rect 254848 495922 254918 495978
rect 254974 495922 255042 495978
rect 255098 495922 255168 495978
rect 254848 495888 255168 495922
rect 285568 496350 285888 496384
rect 285568 496294 285638 496350
rect 285694 496294 285762 496350
rect 285818 496294 285888 496350
rect 285568 496226 285888 496294
rect 285568 496170 285638 496226
rect 285694 496170 285762 496226
rect 285818 496170 285888 496226
rect 285568 496102 285888 496170
rect 285568 496046 285638 496102
rect 285694 496046 285762 496102
rect 285818 496046 285888 496102
rect 285568 495978 285888 496046
rect 285568 495922 285638 495978
rect 285694 495922 285762 495978
rect 285818 495922 285888 495978
rect 285568 495888 285888 495922
rect 316288 496350 316608 496384
rect 316288 496294 316358 496350
rect 316414 496294 316482 496350
rect 316538 496294 316608 496350
rect 316288 496226 316608 496294
rect 316288 496170 316358 496226
rect 316414 496170 316482 496226
rect 316538 496170 316608 496226
rect 316288 496102 316608 496170
rect 316288 496046 316358 496102
rect 316414 496046 316482 496102
rect 316538 496046 316608 496102
rect 316288 495978 316608 496046
rect 316288 495922 316358 495978
rect 316414 495922 316482 495978
rect 316538 495922 316608 495978
rect 316288 495888 316608 495922
rect 347008 496350 347328 496384
rect 347008 496294 347078 496350
rect 347134 496294 347202 496350
rect 347258 496294 347328 496350
rect 347008 496226 347328 496294
rect 347008 496170 347078 496226
rect 347134 496170 347202 496226
rect 347258 496170 347328 496226
rect 347008 496102 347328 496170
rect 347008 496046 347078 496102
rect 347134 496046 347202 496102
rect 347258 496046 347328 496102
rect 347008 495978 347328 496046
rect 347008 495922 347078 495978
rect 347134 495922 347202 495978
rect 347258 495922 347328 495978
rect 347008 495888 347328 495922
rect 377728 496350 378048 496384
rect 377728 496294 377798 496350
rect 377854 496294 377922 496350
rect 377978 496294 378048 496350
rect 377728 496226 378048 496294
rect 377728 496170 377798 496226
rect 377854 496170 377922 496226
rect 377978 496170 378048 496226
rect 377728 496102 378048 496170
rect 377728 496046 377798 496102
rect 377854 496046 377922 496102
rect 377978 496046 378048 496102
rect 377728 495978 378048 496046
rect 377728 495922 377798 495978
rect 377854 495922 377922 495978
rect 377978 495922 378048 495978
rect 377728 495888 378048 495922
rect 408448 496350 408768 496384
rect 408448 496294 408518 496350
rect 408574 496294 408642 496350
rect 408698 496294 408768 496350
rect 408448 496226 408768 496294
rect 408448 496170 408518 496226
rect 408574 496170 408642 496226
rect 408698 496170 408768 496226
rect 408448 496102 408768 496170
rect 408448 496046 408518 496102
rect 408574 496046 408642 496102
rect 408698 496046 408768 496102
rect 408448 495978 408768 496046
rect 408448 495922 408518 495978
rect 408574 495922 408642 495978
rect 408698 495922 408768 495978
rect 408448 495888 408768 495922
rect 439168 496350 439488 496384
rect 439168 496294 439238 496350
rect 439294 496294 439362 496350
rect 439418 496294 439488 496350
rect 439168 496226 439488 496294
rect 439168 496170 439238 496226
rect 439294 496170 439362 496226
rect 439418 496170 439488 496226
rect 439168 496102 439488 496170
rect 439168 496046 439238 496102
rect 439294 496046 439362 496102
rect 439418 496046 439488 496102
rect 439168 495978 439488 496046
rect 439168 495922 439238 495978
rect 439294 495922 439362 495978
rect 439418 495922 439488 495978
rect 439168 495888 439488 495922
rect 469888 496350 470208 496384
rect 469888 496294 469958 496350
rect 470014 496294 470082 496350
rect 470138 496294 470208 496350
rect 469888 496226 470208 496294
rect 469888 496170 469958 496226
rect 470014 496170 470082 496226
rect 470138 496170 470208 496226
rect 469888 496102 470208 496170
rect 469888 496046 469958 496102
rect 470014 496046 470082 496102
rect 470138 496046 470208 496102
rect 469888 495978 470208 496046
rect 469888 495922 469958 495978
rect 470014 495922 470082 495978
rect 470138 495922 470208 495978
rect 469888 495888 470208 495922
rect 500608 496350 500928 496384
rect 500608 496294 500678 496350
rect 500734 496294 500802 496350
rect 500858 496294 500928 496350
rect 500608 496226 500928 496294
rect 500608 496170 500678 496226
rect 500734 496170 500802 496226
rect 500858 496170 500928 496226
rect 500608 496102 500928 496170
rect 500608 496046 500678 496102
rect 500734 496046 500802 496102
rect 500858 496046 500928 496102
rect 500608 495978 500928 496046
rect 500608 495922 500678 495978
rect 500734 495922 500802 495978
rect 500858 495922 500928 495978
rect 500608 495888 500928 495922
rect 24448 490350 24768 490384
rect 24448 490294 24518 490350
rect 24574 490294 24642 490350
rect 24698 490294 24768 490350
rect 24448 490226 24768 490294
rect 24448 490170 24518 490226
rect 24574 490170 24642 490226
rect 24698 490170 24768 490226
rect 24448 490102 24768 490170
rect 24448 490046 24518 490102
rect 24574 490046 24642 490102
rect 24698 490046 24768 490102
rect 24448 489978 24768 490046
rect 24448 489922 24518 489978
rect 24574 489922 24642 489978
rect 24698 489922 24768 489978
rect 24448 489888 24768 489922
rect 55168 490350 55488 490384
rect 55168 490294 55238 490350
rect 55294 490294 55362 490350
rect 55418 490294 55488 490350
rect 55168 490226 55488 490294
rect 55168 490170 55238 490226
rect 55294 490170 55362 490226
rect 55418 490170 55488 490226
rect 55168 490102 55488 490170
rect 55168 490046 55238 490102
rect 55294 490046 55362 490102
rect 55418 490046 55488 490102
rect 55168 489978 55488 490046
rect 55168 489922 55238 489978
rect 55294 489922 55362 489978
rect 55418 489922 55488 489978
rect 55168 489888 55488 489922
rect 85888 490350 86208 490384
rect 85888 490294 85958 490350
rect 86014 490294 86082 490350
rect 86138 490294 86208 490350
rect 85888 490226 86208 490294
rect 85888 490170 85958 490226
rect 86014 490170 86082 490226
rect 86138 490170 86208 490226
rect 85888 490102 86208 490170
rect 85888 490046 85958 490102
rect 86014 490046 86082 490102
rect 86138 490046 86208 490102
rect 85888 489978 86208 490046
rect 85888 489922 85958 489978
rect 86014 489922 86082 489978
rect 86138 489922 86208 489978
rect 85888 489888 86208 489922
rect 116608 490350 116928 490384
rect 116608 490294 116678 490350
rect 116734 490294 116802 490350
rect 116858 490294 116928 490350
rect 116608 490226 116928 490294
rect 116608 490170 116678 490226
rect 116734 490170 116802 490226
rect 116858 490170 116928 490226
rect 116608 490102 116928 490170
rect 116608 490046 116678 490102
rect 116734 490046 116802 490102
rect 116858 490046 116928 490102
rect 116608 489978 116928 490046
rect 116608 489922 116678 489978
rect 116734 489922 116802 489978
rect 116858 489922 116928 489978
rect 116608 489888 116928 489922
rect 147328 490350 147648 490384
rect 147328 490294 147398 490350
rect 147454 490294 147522 490350
rect 147578 490294 147648 490350
rect 147328 490226 147648 490294
rect 147328 490170 147398 490226
rect 147454 490170 147522 490226
rect 147578 490170 147648 490226
rect 147328 490102 147648 490170
rect 147328 490046 147398 490102
rect 147454 490046 147522 490102
rect 147578 490046 147648 490102
rect 147328 489978 147648 490046
rect 147328 489922 147398 489978
rect 147454 489922 147522 489978
rect 147578 489922 147648 489978
rect 147328 489888 147648 489922
rect 178048 490350 178368 490384
rect 178048 490294 178118 490350
rect 178174 490294 178242 490350
rect 178298 490294 178368 490350
rect 178048 490226 178368 490294
rect 178048 490170 178118 490226
rect 178174 490170 178242 490226
rect 178298 490170 178368 490226
rect 178048 490102 178368 490170
rect 178048 490046 178118 490102
rect 178174 490046 178242 490102
rect 178298 490046 178368 490102
rect 178048 489978 178368 490046
rect 178048 489922 178118 489978
rect 178174 489922 178242 489978
rect 178298 489922 178368 489978
rect 178048 489888 178368 489922
rect 208768 490350 209088 490384
rect 208768 490294 208838 490350
rect 208894 490294 208962 490350
rect 209018 490294 209088 490350
rect 208768 490226 209088 490294
rect 208768 490170 208838 490226
rect 208894 490170 208962 490226
rect 209018 490170 209088 490226
rect 208768 490102 209088 490170
rect 208768 490046 208838 490102
rect 208894 490046 208962 490102
rect 209018 490046 209088 490102
rect 208768 489978 209088 490046
rect 208768 489922 208838 489978
rect 208894 489922 208962 489978
rect 209018 489922 209088 489978
rect 208768 489888 209088 489922
rect 239488 490350 239808 490384
rect 239488 490294 239558 490350
rect 239614 490294 239682 490350
rect 239738 490294 239808 490350
rect 239488 490226 239808 490294
rect 239488 490170 239558 490226
rect 239614 490170 239682 490226
rect 239738 490170 239808 490226
rect 239488 490102 239808 490170
rect 239488 490046 239558 490102
rect 239614 490046 239682 490102
rect 239738 490046 239808 490102
rect 239488 489978 239808 490046
rect 239488 489922 239558 489978
rect 239614 489922 239682 489978
rect 239738 489922 239808 489978
rect 239488 489888 239808 489922
rect 270208 490350 270528 490384
rect 270208 490294 270278 490350
rect 270334 490294 270402 490350
rect 270458 490294 270528 490350
rect 270208 490226 270528 490294
rect 270208 490170 270278 490226
rect 270334 490170 270402 490226
rect 270458 490170 270528 490226
rect 270208 490102 270528 490170
rect 270208 490046 270278 490102
rect 270334 490046 270402 490102
rect 270458 490046 270528 490102
rect 270208 489978 270528 490046
rect 270208 489922 270278 489978
rect 270334 489922 270402 489978
rect 270458 489922 270528 489978
rect 270208 489888 270528 489922
rect 300928 490350 301248 490384
rect 300928 490294 300998 490350
rect 301054 490294 301122 490350
rect 301178 490294 301248 490350
rect 300928 490226 301248 490294
rect 300928 490170 300998 490226
rect 301054 490170 301122 490226
rect 301178 490170 301248 490226
rect 300928 490102 301248 490170
rect 300928 490046 300998 490102
rect 301054 490046 301122 490102
rect 301178 490046 301248 490102
rect 300928 489978 301248 490046
rect 300928 489922 300998 489978
rect 301054 489922 301122 489978
rect 301178 489922 301248 489978
rect 300928 489888 301248 489922
rect 331648 490350 331968 490384
rect 331648 490294 331718 490350
rect 331774 490294 331842 490350
rect 331898 490294 331968 490350
rect 331648 490226 331968 490294
rect 331648 490170 331718 490226
rect 331774 490170 331842 490226
rect 331898 490170 331968 490226
rect 331648 490102 331968 490170
rect 331648 490046 331718 490102
rect 331774 490046 331842 490102
rect 331898 490046 331968 490102
rect 331648 489978 331968 490046
rect 331648 489922 331718 489978
rect 331774 489922 331842 489978
rect 331898 489922 331968 489978
rect 331648 489888 331968 489922
rect 362368 490350 362688 490384
rect 362368 490294 362438 490350
rect 362494 490294 362562 490350
rect 362618 490294 362688 490350
rect 362368 490226 362688 490294
rect 362368 490170 362438 490226
rect 362494 490170 362562 490226
rect 362618 490170 362688 490226
rect 362368 490102 362688 490170
rect 362368 490046 362438 490102
rect 362494 490046 362562 490102
rect 362618 490046 362688 490102
rect 362368 489978 362688 490046
rect 362368 489922 362438 489978
rect 362494 489922 362562 489978
rect 362618 489922 362688 489978
rect 362368 489888 362688 489922
rect 393088 490350 393408 490384
rect 393088 490294 393158 490350
rect 393214 490294 393282 490350
rect 393338 490294 393408 490350
rect 393088 490226 393408 490294
rect 393088 490170 393158 490226
rect 393214 490170 393282 490226
rect 393338 490170 393408 490226
rect 393088 490102 393408 490170
rect 393088 490046 393158 490102
rect 393214 490046 393282 490102
rect 393338 490046 393408 490102
rect 393088 489978 393408 490046
rect 393088 489922 393158 489978
rect 393214 489922 393282 489978
rect 393338 489922 393408 489978
rect 393088 489888 393408 489922
rect 423808 490350 424128 490384
rect 423808 490294 423878 490350
rect 423934 490294 424002 490350
rect 424058 490294 424128 490350
rect 423808 490226 424128 490294
rect 423808 490170 423878 490226
rect 423934 490170 424002 490226
rect 424058 490170 424128 490226
rect 423808 490102 424128 490170
rect 423808 490046 423878 490102
rect 423934 490046 424002 490102
rect 424058 490046 424128 490102
rect 423808 489978 424128 490046
rect 423808 489922 423878 489978
rect 423934 489922 424002 489978
rect 424058 489922 424128 489978
rect 423808 489888 424128 489922
rect 454528 490350 454848 490384
rect 454528 490294 454598 490350
rect 454654 490294 454722 490350
rect 454778 490294 454848 490350
rect 454528 490226 454848 490294
rect 454528 490170 454598 490226
rect 454654 490170 454722 490226
rect 454778 490170 454848 490226
rect 454528 490102 454848 490170
rect 454528 490046 454598 490102
rect 454654 490046 454722 490102
rect 454778 490046 454848 490102
rect 454528 489978 454848 490046
rect 454528 489922 454598 489978
rect 454654 489922 454722 489978
rect 454778 489922 454848 489978
rect 454528 489888 454848 489922
rect 485248 490350 485568 490384
rect 485248 490294 485318 490350
rect 485374 490294 485442 490350
rect 485498 490294 485568 490350
rect 485248 490226 485568 490294
rect 485248 490170 485318 490226
rect 485374 490170 485442 490226
rect 485498 490170 485568 490226
rect 485248 490102 485568 490170
rect 485248 490046 485318 490102
rect 485374 490046 485442 490102
rect 485498 490046 485568 490102
rect 485248 489978 485568 490046
rect 485248 489922 485318 489978
rect 485374 489922 485442 489978
rect 485498 489922 485568 489978
rect 485248 489888 485568 489922
rect 515968 490350 516288 490384
rect 515968 490294 516038 490350
rect 516094 490294 516162 490350
rect 516218 490294 516288 490350
rect 515968 490226 516288 490294
rect 515968 490170 516038 490226
rect 516094 490170 516162 490226
rect 516218 490170 516288 490226
rect 515968 490102 516288 490170
rect 515968 490046 516038 490102
rect 516094 490046 516162 490102
rect 516218 490046 516288 490102
rect 515968 489978 516288 490046
rect 515968 489922 516038 489978
rect 516094 489922 516162 489978
rect 516218 489922 516288 489978
rect 515968 489888 516288 489922
rect 525154 490350 525774 507922
rect 525154 490294 525250 490350
rect 525306 490294 525374 490350
rect 525430 490294 525498 490350
rect 525554 490294 525622 490350
rect 525678 490294 525774 490350
rect 525154 490226 525774 490294
rect 525154 490170 525250 490226
rect 525306 490170 525374 490226
rect 525430 490170 525498 490226
rect 525554 490170 525622 490226
rect 525678 490170 525774 490226
rect 525154 490102 525774 490170
rect 525154 490046 525250 490102
rect 525306 490046 525374 490102
rect 525430 490046 525498 490102
rect 525554 490046 525622 490102
rect 525678 490046 525774 490102
rect 525154 489978 525774 490046
rect 525154 489922 525250 489978
rect 525306 489922 525374 489978
rect 525430 489922 525498 489978
rect 525554 489922 525622 489978
rect 525678 489922 525774 489978
rect 6874 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 7494 478350
rect 6874 478226 7494 478294
rect 6874 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 7494 478226
rect 6874 478102 7494 478170
rect 6874 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 7494 478102
rect 6874 477978 7494 478046
rect 6874 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 7494 477978
rect 6874 460350 7494 477922
rect 39808 478350 40128 478384
rect 39808 478294 39878 478350
rect 39934 478294 40002 478350
rect 40058 478294 40128 478350
rect 39808 478226 40128 478294
rect 39808 478170 39878 478226
rect 39934 478170 40002 478226
rect 40058 478170 40128 478226
rect 39808 478102 40128 478170
rect 39808 478046 39878 478102
rect 39934 478046 40002 478102
rect 40058 478046 40128 478102
rect 39808 477978 40128 478046
rect 39808 477922 39878 477978
rect 39934 477922 40002 477978
rect 40058 477922 40128 477978
rect 39808 477888 40128 477922
rect 70528 478350 70848 478384
rect 70528 478294 70598 478350
rect 70654 478294 70722 478350
rect 70778 478294 70848 478350
rect 70528 478226 70848 478294
rect 70528 478170 70598 478226
rect 70654 478170 70722 478226
rect 70778 478170 70848 478226
rect 70528 478102 70848 478170
rect 70528 478046 70598 478102
rect 70654 478046 70722 478102
rect 70778 478046 70848 478102
rect 70528 477978 70848 478046
rect 70528 477922 70598 477978
rect 70654 477922 70722 477978
rect 70778 477922 70848 477978
rect 70528 477888 70848 477922
rect 101248 478350 101568 478384
rect 101248 478294 101318 478350
rect 101374 478294 101442 478350
rect 101498 478294 101568 478350
rect 101248 478226 101568 478294
rect 101248 478170 101318 478226
rect 101374 478170 101442 478226
rect 101498 478170 101568 478226
rect 101248 478102 101568 478170
rect 101248 478046 101318 478102
rect 101374 478046 101442 478102
rect 101498 478046 101568 478102
rect 101248 477978 101568 478046
rect 101248 477922 101318 477978
rect 101374 477922 101442 477978
rect 101498 477922 101568 477978
rect 101248 477888 101568 477922
rect 131968 478350 132288 478384
rect 131968 478294 132038 478350
rect 132094 478294 132162 478350
rect 132218 478294 132288 478350
rect 131968 478226 132288 478294
rect 131968 478170 132038 478226
rect 132094 478170 132162 478226
rect 132218 478170 132288 478226
rect 131968 478102 132288 478170
rect 131968 478046 132038 478102
rect 132094 478046 132162 478102
rect 132218 478046 132288 478102
rect 131968 477978 132288 478046
rect 131968 477922 132038 477978
rect 132094 477922 132162 477978
rect 132218 477922 132288 477978
rect 131968 477888 132288 477922
rect 162688 478350 163008 478384
rect 162688 478294 162758 478350
rect 162814 478294 162882 478350
rect 162938 478294 163008 478350
rect 162688 478226 163008 478294
rect 162688 478170 162758 478226
rect 162814 478170 162882 478226
rect 162938 478170 163008 478226
rect 162688 478102 163008 478170
rect 162688 478046 162758 478102
rect 162814 478046 162882 478102
rect 162938 478046 163008 478102
rect 162688 477978 163008 478046
rect 162688 477922 162758 477978
rect 162814 477922 162882 477978
rect 162938 477922 163008 477978
rect 162688 477888 163008 477922
rect 193408 478350 193728 478384
rect 193408 478294 193478 478350
rect 193534 478294 193602 478350
rect 193658 478294 193728 478350
rect 193408 478226 193728 478294
rect 193408 478170 193478 478226
rect 193534 478170 193602 478226
rect 193658 478170 193728 478226
rect 193408 478102 193728 478170
rect 193408 478046 193478 478102
rect 193534 478046 193602 478102
rect 193658 478046 193728 478102
rect 193408 477978 193728 478046
rect 193408 477922 193478 477978
rect 193534 477922 193602 477978
rect 193658 477922 193728 477978
rect 193408 477888 193728 477922
rect 224128 478350 224448 478384
rect 224128 478294 224198 478350
rect 224254 478294 224322 478350
rect 224378 478294 224448 478350
rect 224128 478226 224448 478294
rect 224128 478170 224198 478226
rect 224254 478170 224322 478226
rect 224378 478170 224448 478226
rect 224128 478102 224448 478170
rect 224128 478046 224198 478102
rect 224254 478046 224322 478102
rect 224378 478046 224448 478102
rect 224128 477978 224448 478046
rect 224128 477922 224198 477978
rect 224254 477922 224322 477978
rect 224378 477922 224448 477978
rect 224128 477888 224448 477922
rect 254848 478350 255168 478384
rect 254848 478294 254918 478350
rect 254974 478294 255042 478350
rect 255098 478294 255168 478350
rect 254848 478226 255168 478294
rect 254848 478170 254918 478226
rect 254974 478170 255042 478226
rect 255098 478170 255168 478226
rect 254848 478102 255168 478170
rect 254848 478046 254918 478102
rect 254974 478046 255042 478102
rect 255098 478046 255168 478102
rect 254848 477978 255168 478046
rect 254848 477922 254918 477978
rect 254974 477922 255042 477978
rect 255098 477922 255168 477978
rect 254848 477888 255168 477922
rect 285568 478350 285888 478384
rect 285568 478294 285638 478350
rect 285694 478294 285762 478350
rect 285818 478294 285888 478350
rect 285568 478226 285888 478294
rect 285568 478170 285638 478226
rect 285694 478170 285762 478226
rect 285818 478170 285888 478226
rect 285568 478102 285888 478170
rect 285568 478046 285638 478102
rect 285694 478046 285762 478102
rect 285818 478046 285888 478102
rect 285568 477978 285888 478046
rect 285568 477922 285638 477978
rect 285694 477922 285762 477978
rect 285818 477922 285888 477978
rect 285568 477888 285888 477922
rect 316288 478350 316608 478384
rect 316288 478294 316358 478350
rect 316414 478294 316482 478350
rect 316538 478294 316608 478350
rect 316288 478226 316608 478294
rect 316288 478170 316358 478226
rect 316414 478170 316482 478226
rect 316538 478170 316608 478226
rect 316288 478102 316608 478170
rect 316288 478046 316358 478102
rect 316414 478046 316482 478102
rect 316538 478046 316608 478102
rect 316288 477978 316608 478046
rect 316288 477922 316358 477978
rect 316414 477922 316482 477978
rect 316538 477922 316608 477978
rect 316288 477888 316608 477922
rect 347008 478350 347328 478384
rect 347008 478294 347078 478350
rect 347134 478294 347202 478350
rect 347258 478294 347328 478350
rect 347008 478226 347328 478294
rect 347008 478170 347078 478226
rect 347134 478170 347202 478226
rect 347258 478170 347328 478226
rect 347008 478102 347328 478170
rect 347008 478046 347078 478102
rect 347134 478046 347202 478102
rect 347258 478046 347328 478102
rect 347008 477978 347328 478046
rect 347008 477922 347078 477978
rect 347134 477922 347202 477978
rect 347258 477922 347328 477978
rect 347008 477888 347328 477922
rect 377728 478350 378048 478384
rect 377728 478294 377798 478350
rect 377854 478294 377922 478350
rect 377978 478294 378048 478350
rect 377728 478226 378048 478294
rect 377728 478170 377798 478226
rect 377854 478170 377922 478226
rect 377978 478170 378048 478226
rect 377728 478102 378048 478170
rect 377728 478046 377798 478102
rect 377854 478046 377922 478102
rect 377978 478046 378048 478102
rect 377728 477978 378048 478046
rect 377728 477922 377798 477978
rect 377854 477922 377922 477978
rect 377978 477922 378048 477978
rect 377728 477888 378048 477922
rect 408448 478350 408768 478384
rect 408448 478294 408518 478350
rect 408574 478294 408642 478350
rect 408698 478294 408768 478350
rect 408448 478226 408768 478294
rect 408448 478170 408518 478226
rect 408574 478170 408642 478226
rect 408698 478170 408768 478226
rect 408448 478102 408768 478170
rect 408448 478046 408518 478102
rect 408574 478046 408642 478102
rect 408698 478046 408768 478102
rect 408448 477978 408768 478046
rect 408448 477922 408518 477978
rect 408574 477922 408642 477978
rect 408698 477922 408768 477978
rect 408448 477888 408768 477922
rect 439168 478350 439488 478384
rect 439168 478294 439238 478350
rect 439294 478294 439362 478350
rect 439418 478294 439488 478350
rect 439168 478226 439488 478294
rect 439168 478170 439238 478226
rect 439294 478170 439362 478226
rect 439418 478170 439488 478226
rect 439168 478102 439488 478170
rect 439168 478046 439238 478102
rect 439294 478046 439362 478102
rect 439418 478046 439488 478102
rect 439168 477978 439488 478046
rect 439168 477922 439238 477978
rect 439294 477922 439362 477978
rect 439418 477922 439488 477978
rect 439168 477888 439488 477922
rect 469888 478350 470208 478384
rect 469888 478294 469958 478350
rect 470014 478294 470082 478350
rect 470138 478294 470208 478350
rect 469888 478226 470208 478294
rect 469888 478170 469958 478226
rect 470014 478170 470082 478226
rect 470138 478170 470208 478226
rect 469888 478102 470208 478170
rect 469888 478046 469958 478102
rect 470014 478046 470082 478102
rect 470138 478046 470208 478102
rect 469888 477978 470208 478046
rect 469888 477922 469958 477978
rect 470014 477922 470082 477978
rect 470138 477922 470208 477978
rect 469888 477888 470208 477922
rect 500608 478350 500928 478384
rect 500608 478294 500678 478350
rect 500734 478294 500802 478350
rect 500858 478294 500928 478350
rect 500608 478226 500928 478294
rect 500608 478170 500678 478226
rect 500734 478170 500802 478226
rect 500858 478170 500928 478226
rect 500608 478102 500928 478170
rect 500608 478046 500678 478102
rect 500734 478046 500802 478102
rect 500858 478046 500928 478102
rect 500608 477978 500928 478046
rect 500608 477922 500678 477978
rect 500734 477922 500802 477978
rect 500858 477922 500928 477978
rect 500608 477888 500928 477922
rect 24448 472350 24768 472384
rect 24448 472294 24518 472350
rect 24574 472294 24642 472350
rect 24698 472294 24768 472350
rect 24448 472226 24768 472294
rect 24448 472170 24518 472226
rect 24574 472170 24642 472226
rect 24698 472170 24768 472226
rect 24448 472102 24768 472170
rect 24448 472046 24518 472102
rect 24574 472046 24642 472102
rect 24698 472046 24768 472102
rect 24448 471978 24768 472046
rect 24448 471922 24518 471978
rect 24574 471922 24642 471978
rect 24698 471922 24768 471978
rect 24448 471888 24768 471922
rect 55168 472350 55488 472384
rect 55168 472294 55238 472350
rect 55294 472294 55362 472350
rect 55418 472294 55488 472350
rect 55168 472226 55488 472294
rect 55168 472170 55238 472226
rect 55294 472170 55362 472226
rect 55418 472170 55488 472226
rect 55168 472102 55488 472170
rect 55168 472046 55238 472102
rect 55294 472046 55362 472102
rect 55418 472046 55488 472102
rect 55168 471978 55488 472046
rect 55168 471922 55238 471978
rect 55294 471922 55362 471978
rect 55418 471922 55488 471978
rect 55168 471888 55488 471922
rect 85888 472350 86208 472384
rect 85888 472294 85958 472350
rect 86014 472294 86082 472350
rect 86138 472294 86208 472350
rect 85888 472226 86208 472294
rect 85888 472170 85958 472226
rect 86014 472170 86082 472226
rect 86138 472170 86208 472226
rect 85888 472102 86208 472170
rect 85888 472046 85958 472102
rect 86014 472046 86082 472102
rect 86138 472046 86208 472102
rect 85888 471978 86208 472046
rect 85888 471922 85958 471978
rect 86014 471922 86082 471978
rect 86138 471922 86208 471978
rect 85888 471888 86208 471922
rect 116608 472350 116928 472384
rect 116608 472294 116678 472350
rect 116734 472294 116802 472350
rect 116858 472294 116928 472350
rect 116608 472226 116928 472294
rect 116608 472170 116678 472226
rect 116734 472170 116802 472226
rect 116858 472170 116928 472226
rect 116608 472102 116928 472170
rect 116608 472046 116678 472102
rect 116734 472046 116802 472102
rect 116858 472046 116928 472102
rect 116608 471978 116928 472046
rect 116608 471922 116678 471978
rect 116734 471922 116802 471978
rect 116858 471922 116928 471978
rect 116608 471888 116928 471922
rect 147328 472350 147648 472384
rect 147328 472294 147398 472350
rect 147454 472294 147522 472350
rect 147578 472294 147648 472350
rect 147328 472226 147648 472294
rect 147328 472170 147398 472226
rect 147454 472170 147522 472226
rect 147578 472170 147648 472226
rect 147328 472102 147648 472170
rect 147328 472046 147398 472102
rect 147454 472046 147522 472102
rect 147578 472046 147648 472102
rect 147328 471978 147648 472046
rect 147328 471922 147398 471978
rect 147454 471922 147522 471978
rect 147578 471922 147648 471978
rect 147328 471888 147648 471922
rect 178048 472350 178368 472384
rect 178048 472294 178118 472350
rect 178174 472294 178242 472350
rect 178298 472294 178368 472350
rect 178048 472226 178368 472294
rect 178048 472170 178118 472226
rect 178174 472170 178242 472226
rect 178298 472170 178368 472226
rect 178048 472102 178368 472170
rect 178048 472046 178118 472102
rect 178174 472046 178242 472102
rect 178298 472046 178368 472102
rect 178048 471978 178368 472046
rect 178048 471922 178118 471978
rect 178174 471922 178242 471978
rect 178298 471922 178368 471978
rect 178048 471888 178368 471922
rect 208768 472350 209088 472384
rect 208768 472294 208838 472350
rect 208894 472294 208962 472350
rect 209018 472294 209088 472350
rect 208768 472226 209088 472294
rect 208768 472170 208838 472226
rect 208894 472170 208962 472226
rect 209018 472170 209088 472226
rect 208768 472102 209088 472170
rect 208768 472046 208838 472102
rect 208894 472046 208962 472102
rect 209018 472046 209088 472102
rect 208768 471978 209088 472046
rect 208768 471922 208838 471978
rect 208894 471922 208962 471978
rect 209018 471922 209088 471978
rect 208768 471888 209088 471922
rect 239488 472350 239808 472384
rect 239488 472294 239558 472350
rect 239614 472294 239682 472350
rect 239738 472294 239808 472350
rect 239488 472226 239808 472294
rect 239488 472170 239558 472226
rect 239614 472170 239682 472226
rect 239738 472170 239808 472226
rect 239488 472102 239808 472170
rect 239488 472046 239558 472102
rect 239614 472046 239682 472102
rect 239738 472046 239808 472102
rect 239488 471978 239808 472046
rect 239488 471922 239558 471978
rect 239614 471922 239682 471978
rect 239738 471922 239808 471978
rect 239488 471888 239808 471922
rect 270208 472350 270528 472384
rect 270208 472294 270278 472350
rect 270334 472294 270402 472350
rect 270458 472294 270528 472350
rect 270208 472226 270528 472294
rect 270208 472170 270278 472226
rect 270334 472170 270402 472226
rect 270458 472170 270528 472226
rect 270208 472102 270528 472170
rect 270208 472046 270278 472102
rect 270334 472046 270402 472102
rect 270458 472046 270528 472102
rect 270208 471978 270528 472046
rect 270208 471922 270278 471978
rect 270334 471922 270402 471978
rect 270458 471922 270528 471978
rect 270208 471888 270528 471922
rect 300928 472350 301248 472384
rect 300928 472294 300998 472350
rect 301054 472294 301122 472350
rect 301178 472294 301248 472350
rect 300928 472226 301248 472294
rect 300928 472170 300998 472226
rect 301054 472170 301122 472226
rect 301178 472170 301248 472226
rect 300928 472102 301248 472170
rect 300928 472046 300998 472102
rect 301054 472046 301122 472102
rect 301178 472046 301248 472102
rect 300928 471978 301248 472046
rect 300928 471922 300998 471978
rect 301054 471922 301122 471978
rect 301178 471922 301248 471978
rect 300928 471888 301248 471922
rect 331648 472350 331968 472384
rect 331648 472294 331718 472350
rect 331774 472294 331842 472350
rect 331898 472294 331968 472350
rect 331648 472226 331968 472294
rect 331648 472170 331718 472226
rect 331774 472170 331842 472226
rect 331898 472170 331968 472226
rect 331648 472102 331968 472170
rect 331648 472046 331718 472102
rect 331774 472046 331842 472102
rect 331898 472046 331968 472102
rect 331648 471978 331968 472046
rect 331648 471922 331718 471978
rect 331774 471922 331842 471978
rect 331898 471922 331968 471978
rect 331648 471888 331968 471922
rect 362368 472350 362688 472384
rect 362368 472294 362438 472350
rect 362494 472294 362562 472350
rect 362618 472294 362688 472350
rect 362368 472226 362688 472294
rect 362368 472170 362438 472226
rect 362494 472170 362562 472226
rect 362618 472170 362688 472226
rect 362368 472102 362688 472170
rect 362368 472046 362438 472102
rect 362494 472046 362562 472102
rect 362618 472046 362688 472102
rect 362368 471978 362688 472046
rect 362368 471922 362438 471978
rect 362494 471922 362562 471978
rect 362618 471922 362688 471978
rect 362368 471888 362688 471922
rect 393088 472350 393408 472384
rect 393088 472294 393158 472350
rect 393214 472294 393282 472350
rect 393338 472294 393408 472350
rect 393088 472226 393408 472294
rect 393088 472170 393158 472226
rect 393214 472170 393282 472226
rect 393338 472170 393408 472226
rect 393088 472102 393408 472170
rect 393088 472046 393158 472102
rect 393214 472046 393282 472102
rect 393338 472046 393408 472102
rect 393088 471978 393408 472046
rect 393088 471922 393158 471978
rect 393214 471922 393282 471978
rect 393338 471922 393408 471978
rect 393088 471888 393408 471922
rect 423808 472350 424128 472384
rect 423808 472294 423878 472350
rect 423934 472294 424002 472350
rect 424058 472294 424128 472350
rect 423808 472226 424128 472294
rect 423808 472170 423878 472226
rect 423934 472170 424002 472226
rect 424058 472170 424128 472226
rect 423808 472102 424128 472170
rect 423808 472046 423878 472102
rect 423934 472046 424002 472102
rect 424058 472046 424128 472102
rect 423808 471978 424128 472046
rect 423808 471922 423878 471978
rect 423934 471922 424002 471978
rect 424058 471922 424128 471978
rect 423808 471888 424128 471922
rect 454528 472350 454848 472384
rect 454528 472294 454598 472350
rect 454654 472294 454722 472350
rect 454778 472294 454848 472350
rect 454528 472226 454848 472294
rect 454528 472170 454598 472226
rect 454654 472170 454722 472226
rect 454778 472170 454848 472226
rect 454528 472102 454848 472170
rect 454528 472046 454598 472102
rect 454654 472046 454722 472102
rect 454778 472046 454848 472102
rect 454528 471978 454848 472046
rect 454528 471922 454598 471978
rect 454654 471922 454722 471978
rect 454778 471922 454848 471978
rect 454528 471888 454848 471922
rect 485248 472350 485568 472384
rect 485248 472294 485318 472350
rect 485374 472294 485442 472350
rect 485498 472294 485568 472350
rect 485248 472226 485568 472294
rect 485248 472170 485318 472226
rect 485374 472170 485442 472226
rect 485498 472170 485568 472226
rect 485248 472102 485568 472170
rect 485248 472046 485318 472102
rect 485374 472046 485442 472102
rect 485498 472046 485568 472102
rect 485248 471978 485568 472046
rect 485248 471922 485318 471978
rect 485374 471922 485442 471978
rect 485498 471922 485568 471978
rect 485248 471888 485568 471922
rect 515968 472350 516288 472384
rect 515968 472294 516038 472350
rect 516094 472294 516162 472350
rect 516218 472294 516288 472350
rect 515968 472226 516288 472294
rect 515968 472170 516038 472226
rect 516094 472170 516162 472226
rect 516218 472170 516288 472226
rect 515968 472102 516288 472170
rect 515968 472046 516038 472102
rect 516094 472046 516162 472102
rect 516218 472046 516288 472102
rect 515968 471978 516288 472046
rect 515968 471922 516038 471978
rect 516094 471922 516162 471978
rect 516218 471922 516288 471978
rect 515968 471888 516288 471922
rect 525154 472350 525774 489922
rect 525154 472294 525250 472350
rect 525306 472294 525374 472350
rect 525430 472294 525498 472350
rect 525554 472294 525622 472350
rect 525678 472294 525774 472350
rect 525154 472226 525774 472294
rect 525154 472170 525250 472226
rect 525306 472170 525374 472226
rect 525430 472170 525498 472226
rect 525554 472170 525622 472226
rect 525678 472170 525774 472226
rect 525154 472102 525774 472170
rect 525154 472046 525250 472102
rect 525306 472046 525374 472102
rect 525430 472046 525498 472102
rect 525554 472046 525622 472102
rect 525678 472046 525774 472102
rect 525154 471978 525774 472046
rect 525154 471922 525250 471978
rect 525306 471922 525374 471978
rect 525430 471922 525498 471978
rect 525554 471922 525622 471978
rect 525678 471922 525774 471978
rect 6874 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 7494 460350
rect 6874 460226 7494 460294
rect 6874 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 7494 460226
rect 6874 460102 7494 460170
rect 6874 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 7494 460102
rect 6874 459978 7494 460046
rect 6874 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 7494 459978
rect 6874 442350 7494 459922
rect 39808 460350 40128 460384
rect 39808 460294 39878 460350
rect 39934 460294 40002 460350
rect 40058 460294 40128 460350
rect 39808 460226 40128 460294
rect 39808 460170 39878 460226
rect 39934 460170 40002 460226
rect 40058 460170 40128 460226
rect 39808 460102 40128 460170
rect 39808 460046 39878 460102
rect 39934 460046 40002 460102
rect 40058 460046 40128 460102
rect 39808 459978 40128 460046
rect 39808 459922 39878 459978
rect 39934 459922 40002 459978
rect 40058 459922 40128 459978
rect 39808 459888 40128 459922
rect 70528 460350 70848 460384
rect 70528 460294 70598 460350
rect 70654 460294 70722 460350
rect 70778 460294 70848 460350
rect 70528 460226 70848 460294
rect 70528 460170 70598 460226
rect 70654 460170 70722 460226
rect 70778 460170 70848 460226
rect 70528 460102 70848 460170
rect 70528 460046 70598 460102
rect 70654 460046 70722 460102
rect 70778 460046 70848 460102
rect 70528 459978 70848 460046
rect 70528 459922 70598 459978
rect 70654 459922 70722 459978
rect 70778 459922 70848 459978
rect 70528 459888 70848 459922
rect 101248 460350 101568 460384
rect 101248 460294 101318 460350
rect 101374 460294 101442 460350
rect 101498 460294 101568 460350
rect 101248 460226 101568 460294
rect 101248 460170 101318 460226
rect 101374 460170 101442 460226
rect 101498 460170 101568 460226
rect 101248 460102 101568 460170
rect 101248 460046 101318 460102
rect 101374 460046 101442 460102
rect 101498 460046 101568 460102
rect 101248 459978 101568 460046
rect 101248 459922 101318 459978
rect 101374 459922 101442 459978
rect 101498 459922 101568 459978
rect 101248 459888 101568 459922
rect 131968 460350 132288 460384
rect 131968 460294 132038 460350
rect 132094 460294 132162 460350
rect 132218 460294 132288 460350
rect 131968 460226 132288 460294
rect 131968 460170 132038 460226
rect 132094 460170 132162 460226
rect 132218 460170 132288 460226
rect 131968 460102 132288 460170
rect 131968 460046 132038 460102
rect 132094 460046 132162 460102
rect 132218 460046 132288 460102
rect 131968 459978 132288 460046
rect 131968 459922 132038 459978
rect 132094 459922 132162 459978
rect 132218 459922 132288 459978
rect 131968 459888 132288 459922
rect 162688 460350 163008 460384
rect 162688 460294 162758 460350
rect 162814 460294 162882 460350
rect 162938 460294 163008 460350
rect 162688 460226 163008 460294
rect 162688 460170 162758 460226
rect 162814 460170 162882 460226
rect 162938 460170 163008 460226
rect 162688 460102 163008 460170
rect 162688 460046 162758 460102
rect 162814 460046 162882 460102
rect 162938 460046 163008 460102
rect 162688 459978 163008 460046
rect 162688 459922 162758 459978
rect 162814 459922 162882 459978
rect 162938 459922 163008 459978
rect 162688 459888 163008 459922
rect 193408 460350 193728 460384
rect 193408 460294 193478 460350
rect 193534 460294 193602 460350
rect 193658 460294 193728 460350
rect 193408 460226 193728 460294
rect 193408 460170 193478 460226
rect 193534 460170 193602 460226
rect 193658 460170 193728 460226
rect 193408 460102 193728 460170
rect 193408 460046 193478 460102
rect 193534 460046 193602 460102
rect 193658 460046 193728 460102
rect 193408 459978 193728 460046
rect 193408 459922 193478 459978
rect 193534 459922 193602 459978
rect 193658 459922 193728 459978
rect 193408 459888 193728 459922
rect 224128 460350 224448 460384
rect 224128 460294 224198 460350
rect 224254 460294 224322 460350
rect 224378 460294 224448 460350
rect 224128 460226 224448 460294
rect 224128 460170 224198 460226
rect 224254 460170 224322 460226
rect 224378 460170 224448 460226
rect 224128 460102 224448 460170
rect 224128 460046 224198 460102
rect 224254 460046 224322 460102
rect 224378 460046 224448 460102
rect 224128 459978 224448 460046
rect 224128 459922 224198 459978
rect 224254 459922 224322 459978
rect 224378 459922 224448 459978
rect 224128 459888 224448 459922
rect 254848 460350 255168 460384
rect 254848 460294 254918 460350
rect 254974 460294 255042 460350
rect 255098 460294 255168 460350
rect 254848 460226 255168 460294
rect 254848 460170 254918 460226
rect 254974 460170 255042 460226
rect 255098 460170 255168 460226
rect 254848 460102 255168 460170
rect 254848 460046 254918 460102
rect 254974 460046 255042 460102
rect 255098 460046 255168 460102
rect 254848 459978 255168 460046
rect 254848 459922 254918 459978
rect 254974 459922 255042 459978
rect 255098 459922 255168 459978
rect 254848 459888 255168 459922
rect 285568 460350 285888 460384
rect 285568 460294 285638 460350
rect 285694 460294 285762 460350
rect 285818 460294 285888 460350
rect 285568 460226 285888 460294
rect 285568 460170 285638 460226
rect 285694 460170 285762 460226
rect 285818 460170 285888 460226
rect 285568 460102 285888 460170
rect 285568 460046 285638 460102
rect 285694 460046 285762 460102
rect 285818 460046 285888 460102
rect 285568 459978 285888 460046
rect 285568 459922 285638 459978
rect 285694 459922 285762 459978
rect 285818 459922 285888 459978
rect 285568 459888 285888 459922
rect 316288 460350 316608 460384
rect 316288 460294 316358 460350
rect 316414 460294 316482 460350
rect 316538 460294 316608 460350
rect 316288 460226 316608 460294
rect 316288 460170 316358 460226
rect 316414 460170 316482 460226
rect 316538 460170 316608 460226
rect 316288 460102 316608 460170
rect 316288 460046 316358 460102
rect 316414 460046 316482 460102
rect 316538 460046 316608 460102
rect 316288 459978 316608 460046
rect 316288 459922 316358 459978
rect 316414 459922 316482 459978
rect 316538 459922 316608 459978
rect 316288 459888 316608 459922
rect 347008 460350 347328 460384
rect 347008 460294 347078 460350
rect 347134 460294 347202 460350
rect 347258 460294 347328 460350
rect 347008 460226 347328 460294
rect 347008 460170 347078 460226
rect 347134 460170 347202 460226
rect 347258 460170 347328 460226
rect 347008 460102 347328 460170
rect 347008 460046 347078 460102
rect 347134 460046 347202 460102
rect 347258 460046 347328 460102
rect 347008 459978 347328 460046
rect 347008 459922 347078 459978
rect 347134 459922 347202 459978
rect 347258 459922 347328 459978
rect 347008 459888 347328 459922
rect 377728 460350 378048 460384
rect 377728 460294 377798 460350
rect 377854 460294 377922 460350
rect 377978 460294 378048 460350
rect 377728 460226 378048 460294
rect 377728 460170 377798 460226
rect 377854 460170 377922 460226
rect 377978 460170 378048 460226
rect 377728 460102 378048 460170
rect 377728 460046 377798 460102
rect 377854 460046 377922 460102
rect 377978 460046 378048 460102
rect 377728 459978 378048 460046
rect 377728 459922 377798 459978
rect 377854 459922 377922 459978
rect 377978 459922 378048 459978
rect 377728 459888 378048 459922
rect 408448 460350 408768 460384
rect 408448 460294 408518 460350
rect 408574 460294 408642 460350
rect 408698 460294 408768 460350
rect 408448 460226 408768 460294
rect 408448 460170 408518 460226
rect 408574 460170 408642 460226
rect 408698 460170 408768 460226
rect 408448 460102 408768 460170
rect 408448 460046 408518 460102
rect 408574 460046 408642 460102
rect 408698 460046 408768 460102
rect 408448 459978 408768 460046
rect 408448 459922 408518 459978
rect 408574 459922 408642 459978
rect 408698 459922 408768 459978
rect 408448 459888 408768 459922
rect 439168 460350 439488 460384
rect 439168 460294 439238 460350
rect 439294 460294 439362 460350
rect 439418 460294 439488 460350
rect 439168 460226 439488 460294
rect 439168 460170 439238 460226
rect 439294 460170 439362 460226
rect 439418 460170 439488 460226
rect 439168 460102 439488 460170
rect 439168 460046 439238 460102
rect 439294 460046 439362 460102
rect 439418 460046 439488 460102
rect 439168 459978 439488 460046
rect 439168 459922 439238 459978
rect 439294 459922 439362 459978
rect 439418 459922 439488 459978
rect 439168 459888 439488 459922
rect 469888 460350 470208 460384
rect 469888 460294 469958 460350
rect 470014 460294 470082 460350
rect 470138 460294 470208 460350
rect 469888 460226 470208 460294
rect 469888 460170 469958 460226
rect 470014 460170 470082 460226
rect 470138 460170 470208 460226
rect 469888 460102 470208 460170
rect 469888 460046 469958 460102
rect 470014 460046 470082 460102
rect 470138 460046 470208 460102
rect 469888 459978 470208 460046
rect 469888 459922 469958 459978
rect 470014 459922 470082 459978
rect 470138 459922 470208 459978
rect 469888 459888 470208 459922
rect 500608 460350 500928 460384
rect 500608 460294 500678 460350
rect 500734 460294 500802 460350
rect 500858 460294 500928 460350
rect 500608 460226 500928 460294
rect 500608 460170 500678 460226
rect 500734 460170 500802 460226
rect 500858 460170 500928 460226
rect 500608 460102 500928 460170
rect 500608 460046 500678 460102
rect 500734 460046 500802 460102
rect 500858 460046 500928 460102
rect 500608 459978 500928 460046
rect 500608 459922 500678 459978
rect 500734 459922 500802 459978
rect 500858 459922 500928 459978
rect 500608 459888 500928 459922
rect 24448 454350 24768 454384
rect 24448 454294 24518 454350
rect 24574 454294 24642 454350
rect 24698 454294 24768 454350
rect 24448 454226 24768 454294
rect 24448 454170 24518 454226
rect 24574 454170 24642 454226
rect 24698 454170 24768 454226
rect 24448 454102 24768 454170
rect 24448 454046 24518 454102
rect 24574 454046 24642 454102
rect 24698 454046 24768 454102
rect 24448 453978 24768 454046
rect 24448 453922 24518 453978
rect 24574 453922 24642 453978
rect 24698 453922 24768 453978
rect 24448 453888 24768 453922
rect 55168 454350 55488 454384
rect 55168 454294 55238 454350
rect 55294 454294 55362 454350
rect 55418 454294 55488 454350
rect 55168 454226 55488 454294
rect 55168 454170 55238 454226
rect 55294 454170 55362 454226
rect 55418 454170 55488 454226
rect 55168 454102 55488 454170
rect 55168 454046 55238 454102
rect 55294 454046 55362 454102
rect 55418 454046 55488 454102
rect 55168 453978 55488 454046
rect 55168 453922 55238 453978
rect 55294 453922 55362 453978
rect 55418 453922 55488 453978
rect 55168 453888 55488 453922
rect 85888 454350 86208 454384
rect 85888 454294 85958 454350
rect 86014 454294 86082 454350
rect 86138 454294 86208 454350
rect 85888 454226 86208 454294
rect 85888 454170 85958 454226
rect 86014 454170 86082 454226
rect 86138 454170 86208 454226
rect 85888 454102 86208 454170
rect 85888 454046 85958 454102
rect 86014 454046 86082 454102
rect 86138 454046 86208 454102
rect 85888 453978 86208 454046
rect 85888 453922 85958 453978
rect 86014 453922 86082 453978
rect 86138 453922 86208 453978
rect 85888 453888 86208 453922
rect 116608 454350 116928 454384
rect 116608 454294 116678 454350
rect 116734 454294 116802 454350
rect 116858 454294 116928 454350
rect 116608 454226 116928 454294
rect 116608 454170 116678 454226
rect 116734 454170 116802 454226
rect 116858 454170 116928 454226
rect 116608 454102 116928 454170
rect 116608 454046 116678 454102
rect 116734 454046 116802 454102
rect 116858 454046 116928 454102
rect 116608 453978 116928 454046
rect 116608 453922 116678 453978
rect 116734 453922 116802 453978
rect 116858 453922 116928 453978
rect 116608 453888 116928 453922
rect 147328 454350 147648 454384
rect 147328 454294 147398 454350
rect 147454 454294 147522 454350
rect 147578 454294 147648 454350
rect 147328 454226 147648 454294
rect 147328 454170 147398 454226
rect 147454 454170 147522 454226
rect 147578 454170 147648 454226
rect 147328 454102 147648 454170
rect 147328 454046 147398 454102
rect 147454 454046 147522 454102
rect 147578 454046 147648 454102
rect 147328 453978 147648 454046
rect 147328 453922 147398 453978
rect 147454 453922 147522 453978
rect 147578 453922 147648 453978
rect 147328 453888 147648 453922
rect 178048 454350 178368 454384
rect 178048 454294 178118 454350
rect 178174 454294 178242 454350
rect 178298 454294 178368 454350
rect 178048 454226 178368 454294
rect 178048 454170 178118 454226
rect 178174 454170 178242 454226
rect 178298 454170 178368 454226
rect 178048 454102 178368 454170
rect 178048 454046 178118 454102
rect 178174 454046 178242 454102
rect 178298 454046 178368 454102
rect 178048 453978 178368 454046
rect 178048 453922 178118 453978
rect 178174 453922 178242 453978
rect 178298 453922 178368 453978
rect 178048 453888 178368 453922
rect 208768 454350 209088 454384
rect 208768 454294 208838 454350
rect 208894 454294 208962 454350
rect 209018 454294 209088 454350
rect 208768 454226 209088 454294
rect 208768 454170 208838 454226
rect 208894 454170 208962 454226
rect 209018 454170 209088 454226
rect 208768 454102 209088 454170
rect 208768 454046 208838 454102
rect 208894 454046 208962 454102
rect 209018 454046 209088 454102
rect 208768 453978 209088 454046
rect 208768 453922 208838 453978
rect 208894 453922 208962 453978
rect 209018 453922 209088 453978
rect 208768 453888 209088 453922
rect 239488 454350 239808 454384
rect 239488 454294 239558 454350
rect 239614 454294 239682 454350
rect 239738 454294 239808 454350
rect 239488 454226 239808 454294
rect 239488 454170 239558 454226
rect 239614 454170 239682 454226
rect 239738 454170 239808 454226
rect 239488 454102 239808 454170
rect 239488 454046 239558 454102
rect 239614 454046 239682 454102
rect 239738 454046 239808 454102
rect 239488 453978 239808 454046
rect 239488 453922 239558 453978
rect 239614 453922 239682 453978
rect 239738 453922 239808 453978
rect 239488 453888 239808 453922
rect 270208 454350 270528 454384
rect 270208 454294 270278 454350
rect 270334 454294 270402 454350
rect 270458 454294 270528 454350
rect 270208 454226 270528 454294
rect 270208 454170 270278 454226
rect 270334 454170 270402 454226
rect 270458 454170 270528 454226
rect 270208 454102 270528 454170
rect 270208 454046 270278 454102
rect 270334 454046 270402 454102
rect 270458 454046 270528 454102
rect 270208 453978 270528 454046
rect 270208 453922 270278 453978
rect 270334 453922 270402 453978
rect 270458 453922 270528 453978
rect 270208 453888 270528 453922
rect 300928 454350 301248 454384
rect 300928 454294 300998 454350
rect 301054 454294 301122 454350
rect 301178 454294 301248 454350
rect 300928 454226 301248 454294
rect 300928 454170 300998 454226
rect 301054 454170 301122 454226
rect 301178 454170 301248 454226
rect 300928 454102 301248 454170
rect 300928 454046 300998 454102
rect 301054 454046 301122 454102
rect 301178 454046 301248 454102
rect 300928 453978 301248 454046
rect 300928 453922 300998 453978
rect 301054 453922 301122 453978
rect 301178 453922 301248 453978
rect 300928 453888 301248 453922
rect 331648 454350 331968 454384
rect 331648 454294 331718 454350
rect 331774 454294 331842 454350
rect 331898 454294 331968 454350
rect 331648 454226 331968 454294
rect 331648 454170 331718 454226
rect 331774 454170 331842 454226
rect 331898 454170 331968 454226
rect 331648 454102 331968 454170
rect 331648 454046 331718 454102
rect 331774 454046 331842 454102
rect 331898 454046 331968 454102
rect 331648 453978 331968 454046
rect 331648 453922 331718 453978
rect 331774 453922 331842 453978
rect 331898 453922 331968 453978
rect 331648 453888 331968 453922
rect 362368 454350 362688 454384
rect 362368 454294 362438 454350
rect 362494 454294 362562 454350
rect 362618 454294 362688 454350
rect 362368 454226 362688 454294
rect 362368 454170 362438 454226
rect 362494 454170 362562 454226
rect 362618 454170 362688 454226
rect 362368 454102 362688 454170
rect 362368 454046 362438 454102
rect 362494 454046 362562 454102
rect 362618 454046 362688 454102
rect 362368 453978 362688 454046
rect 362368 453922 362438 453978
rect 362494 453922 362562 453978
rect 362618 453922 362688 453978
rect 362368 453888 362688 453922
rect 393088 454350 393408 454384
rect 393088 454294 393158 454350
rect 393214 454294 393282 454350
rect 393338 454294 393408 454350
rect 393088 454226 393408 454294
rect 393088 454170 393158 454226
rect 393214 454170 393282 454226
rect 393338 454170 393408 454226
rect 393088 454102 393408 454170
rect 393088 454046 393158 454102
rect 393214 454046 393282 454102
rect 393338 454046 393408 454102
rect 393088 453978 393408 454046
rect 393088 453922 393158 453978
rect 393214 453922 393282 453978
rect 393338 453922 393408 453978
rect 393088 453888 393408 453922
rect 423808 454350 424128 454384
rect 423808 454294 423878 454350
rect 423934 454294 424002 454350
rect 424058 454294 424128 454350
rect 423808 454226 424128 454294
rect 423808 454170 423878 454226
rect 423934 454170 424002 454226
rect 424058 454170 424128 454226
rect 423808 454102 424128 454170
rect 423808 454046 423878 454102
rect 423934 454046 424002 454102
rect 424058 454046 424128 454102
rect 423808 453978 424128 454046
rect 423808 453922 423878 453978
rect 423934 453922 424002 453978
rect 424058 453922 424128 453978
rect 423808 453888 424128 453922
rect 454528 454350 454848 454384
rect 454528 454294 454598 454350
rect 454654 454294 454722 454350
rect 454778 454294 454848 454350
rect 454528 454226 454848 454294
rect 454528 454170 454598 454226
rect 454654 454170 454722 454226
rect 454778 454170 454848 454226
rect 454528 454102 454848 454170
rect 454528 454046 454598 454102
rect 454654 454046 454722 454102
rect 454778 454046 454848 454102
rect 454528 453978 454848 454046
rect 454528 453922 454598 453978
rect 454654 453922 454722 453978
rect 454778 453922 454848 453978
rect 454528 453888 454848 453922
rect 485248 454350 485568 454384
rect 485248 454294 485318 454350
rect 485374 454294 485442 454350
rect 485498 454294 485568 454350
rect 485248 454226 485568 454294
rect 485248 454170 485318 454226
rect 485374 454170 485442 454226
rect 485498 454170 485568 454226
rect 485248 454102 485568 454170
rect 485248 454046 485318 454102
rect 485374 454046 485442 454102
rect 485498 454046 485568 454102
rect 485248 453978 485568 454046
rect 485248 453922 485318 453978
rect 485374 453922 485442 453978
rect 485498 453922 485568 453978
rect 485248 453888 485568 453922
rect 515968 454350 516288 454384
rect 515968 454294 516038 454350
rect 516094 454294 516162 454350
rect 516218 454294 516288 454350
rect 515968 454226 516288 454294
rect 515968 454170 516038 454226
rect 516094 454170 516162 454226
rect 516218 454170 516288 454226
rect 515968 454102 516288 454170
rect 515968 454046 516038 454102
rect 516094 454046 516162 454102
rect 516218 454046 516288 454102
rect 515968 453978 516288 454046
rect 515968 453922 516038 453978
rect 516094 453922 516162 453978
rect 516218 453922 516288 453978
rect 515968 453888 516288 453922
rect 525154 454350 525774 471922
rect 525154 454294 525250 454350
rect 525306 454294 525374 454350
rect 525430 454294 525498 454350
rect 525554 454294 525622 454350
rect 525678 454294 525774 454350
rect 525154 454226 525774 454294
rect 525154 454170 525250 454226
rect 525306 454170 525374 454226
rect 525430 454170 525498 454226
rect 525554 454170 525622 454226
rect 525678 454170 525774 454226
rect 525154 454102 525774 454170
rect 525154 454046 525250 454102
rect 525306 454046 525374 454102
rect 525430 454046 525498 454102
rect 525554 454046 525622 454102
rect 525678 454046 525774 454102
rect 525154 453978 525774 454046
rect 525154 453922 525250 453978
rect 525306 453922 525374 453978
rect 525430 453922 525498 453978
rect 525554 453922 525622 453978
rect 525678 453922 525774 453978
rect 6874 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 7494 442350
rect 6874 442226 7494 442294
rect 6874 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 7494 442226
rect 6874 442102 7494 442170
rect 6874 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 7494 442102
rect 6874 441978 7494 442046
rect 6874 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 7494 441978
rect 6874 424350 7494 441922
rect 39808 442350 40128 442384
rect 39808 442294 39878 442350
rect 39934 442294 40002 442350
rect 40058 442294 40128 442350
rect 39808 442226 40128 442294
rect 39808 442170 39878 442226
rect 39934 442170 40002 442226
rect 40058 442170 40128 442226
rect 39808 442102 40128 442170
rect 39808 442046 39878 442102
rect 39934 442046 40002 442102
rect 40058 442046 40128 442102
rect 39808 441978 40128 442046
rect 39808 441922 39878 441978
rect 39934 441922 40002 441978
rect 40058 441922 40128 441978
rect 39808 441888 40128 441922
rect 70528 442350 70848 442384
rect 70528 442294 70598 442350
rect 70654 442294 70722 442350
rect 70778 442294 70848 442350
rect 70528 442226 70848 442294
rect 70528 442170 70598 442226
rect 70654 442170 70722 442226
rect 70778 442170 70848 442226
rect 70528 442102 70848 442170
rect 70528 442046 70598 442102
rect 70654 442046 70722 442102
rect 70778 442046 70848 442102
rect 70528 441978 70848 442046
rect 70528 441922 70598 441978
rect 70654 441922 70722 441978
rect 70778 441922 70848 441978
rect 70528 441888 70848 441922
rect 101248 442350 101568 442384
rect 101248 442294 101318 442350
rect 101374 442294 101442 442350
rect 101498 442294 101568 442350
rect 101248 442226 101568 442294
rect 101248 442170 101318 442226
rect 101374 442170 101442 442226
rect 101498 442170 101568 442226
rect 101248 442102 101568 442170
rect 101248 442046 101318 442102
rect 101374 442046 101442 442102
rect 101498 442046 101568 442102
rect 101248 441978 101568 442046
rect 101248 441922 101318 441978
rect 101374 441922 101442 441978
rect 101498 441922 101568 441978
rect 101248 441888 101568 441922
rect 131968 442350 132288 442384
rect 131968 442294 132038 442350
rect 132094 442294 132162 442350
rect 132218 442294 132288 442350
rect 131968 442226 132288 442294
rect 131968 442170 132038 442226
rect 132094 442170 132162 442226
rect 132218 442170 132288 442226
rect 131968 442102 132288 442170
rect 131968 442046 132038 442102
rect 132094 442046 132162 442102
rect 132218 442046 132288 442102
rect 131968 441978 132288 442046
rect 131968 441922 132038 441978
rect 132094 441922 132162 441978
rect 132218 441922 132288 441978
rect 131968 441888 132288 441922
rect 162688 442350 163008 442384
rect 162688 442294 162758 442350
rect 162814 442294 162882 442350
rect 162938 442294 163008 442350
rect 162688 442226 163008 442294
rect 162688 442170 162758 442226
rect 162814 442170 162882 442226
rect 162938 442170 163008 442226
rect 162688 442102 163008 442170
rect 162688 442046 162758 442102
rect 162814 442046 162882 442102
rect 162938 442046 163008 442102
rect 162688 441978 163008 442046
rect 162688 441922 162758 441978
rect 162814 441922 162882 441978
rect 162938 441922 163008 441978
rect 162688 441888 163008 441922
rect 193408 442350 193728 442384
rect 193408 442294 193478 442350
rect 193534 442294 193602 442350
rect 193658 442294 193728 442350
rect 193408 442226 193728 442294
rect 193408 442170 193478 442226
rect 193534 442170 193602 442226
rect 193658 442170 193728 442226
rect 193408 442102 193728 442170
rect 193408 442046 193478 442102
rect 193534 442046 193602 442102
rect 193658 442046 193728 442102
rect 193408 441978 193728 442046
rect 193408 441922 193478 441978
rect 193534 441922 193602 441978
rect 193658 441922 193728 441978
rect 193408 441888 193728 441922
rect 224128 442350 224448 442384
rect 224128 442294 224198 442350
rect 224254 442294 224322 442350
rect 224378 442294 224448 442350
rect 224128 442226 224448 442294
rect 224128 442170 224198 442226
rect 224254 442170 224322 442226
rect 224378 442170 224448 442226
rect 224128 442102 224448 442170
rect 224128 442046 224198 442102
rect 224254 442046 224322 442102
rect 224378 442046 224448 442102
rect 224128 441978 224448 442046
rect 224128 441922 224198 441978
rect 224254 441922 224322 441978
rect 224378 441922 224448 441978
rect 224128 441888 224448 441922
rect 254848 442350 255168 442384
rect 254848 442294 254918 442350
rect 254974 442294 255042 442350
rect 255098 442294 255168 442350
rect 254848 442226 255168 442294
rect 254848 442170 254918 442226
rect 254974 442170 255042 442226
rect 255098 442170 255168 442226
rect 254848 442102 255168 442170
rect 254848 442046 254918 442102
rect 254974 442046 255042 442102
rect 255098 442046 255168 442102
rect 254848 441978 255168 442046
rect 254848 441922 254918 441978
rect 254974 441922 255042 441978
rect 255098 441922 255168 441978
rect 254848 441888 255168 441922
rect 285568 442350 285888 442384
rect 285568 442294 285638 442350
rect 285694 442294 285762 442350
rect 285818 442294 285888 442350
rect 285568 442226 285888 442294
rect 285568 442170 285638 442226
rect 285694 442170 285762 442226
rect 285818 442170 285888 442226
rect 285568 442102 285888 442170
rect 285568 442046 285638 442102
rect 285694 442046 285762 442102
rect 285818 442046 285888 442102
rect 285568 441978 285888 442046
rect 285568 441922 285638 441978
rect 285694 441922 285762 441978
rect 285818 441922 285888 441978
rect 285568 441888 285888 441922
rect 316288 442350 316608 442384
rect 316288 442294 316358 442350
rect 316414 442294 316482 442350
rect 316538 442294 316608 442350
rect 316288 442226 316608 442294
rect 316288 442170 316358 442226
rect 316414 442170 316482 442226
rect 316538 442170 316608 442226
rect 316288 442102 316608 442170
rect 316288 442046 316358 442102
rect 316414 442046 316482 442102
rect 316538 442046 316608 442102
rect 316288 441978 316608 442046
rect 316288 441922 316358 441978
rect 316414 441922 316482 441978
rect 316538 441922 316608 441978
rect 316288 441888 316608 441922
rect 347008 442350 347328 442384
rect 347008 442294 347078 442350
rect 347134 442294 347202 442350
rect 347258 442294 347328 442350
rect 347008 442226 347328 442294
rect 347008 442170 347078 442226
rect 347134 442170 347202 442226
rect 347258 442170 347328 442226
rect 347008 442102 347328 442170
rect 347008 442046 347078 442102
rect 347134 442046 347202 442102
rect 347258 442046 347328 442102
rect 347008 441978 347328 442046
rect 347008 441922 347078 441978
rect 347134 441922 347202 441978
rect 347258 441922 347328 441978
rect 347008 441888 347328 441922
rect 377728 442350 378048 442384
rect 377728 442294 377798 442350
rect 377854 442294 377922 442350
rect 377978 442294 378048 442350
rect 377728 442226 378048 442294
rect 377728 442170 377798 442226
rect 377854 442170 377922 442226
rect 377978 442170 378048 442226
rect 377728 442102 378048 442170
rect 377728 442046 377798 442102
rect 377854 442046 377922 442102
rect 377978 442046 378048 442102
rect 377728 441978 378048 442046
rect 377728 441922 377798 441978
rect 377854 441922 377922 441978
rect 377978 441922 378048 441978
rect 377728 441888 378048 441922
rect 408448 442350 408768 442384
rect 408448 442294 408518 442350
rect 408574 442294 408642 442350
rect 408698 442294 408768 442350
rect 408448 442226 408768 442294
rect 408448 442170 408518 442226
rect 408574 442170 408642 442226
rect 408698 442170 408768 442226
rect 408448 442102 408768 442170
rect 408448 442046 408518 442102
rect 408574 442046 408642 442102
rect 408698 442046 408768 442102
rect 408448 441978 408768 442046
rect 408448 441922 408518 441978
rect 408574 441922 408642 441978
rect 408698 441922 408768 441978
rect 408448 441888 408768 441922
rect 439168 442350 439488 442384
rect 439168 442294 439238 442350
rect 439294 442294 439362 442350
rect 439418 442294 439488 442350
rect 439168 442226 439488 442294
rect 439168 442170 439238 442226
rect 439294 442170 439362 442226
rect 439418 442170 439488 442226
rect 439168 442102 439488 442170
rect 439168 442046 439238 442102
rect 439294 442046 439362 442102
rect 439418 442046 439488 442102
rect 439168 441978 439488 442046
rect 439168 441922 439238 441978
rect 439294 441922 439362 441978
rect 439418 441922 439488 441978
rect 439168 441888 439488 441922
rect 469888 442350 470208 442384
rect 469888 442294 469958 442350
rect 470014 442294 470082 442350
rect 470138 442294 470208 442350
rect 469888 442226 470208 442294
rect 469888 442170 469958 442226
rect 470014 442170 470082 442226
rect 470138 442170 470208 442226
rect 469888 442102 470208 442170
rect 469888 442046 469958 442102
rect 470014 442046 470082 442102
rect 470138 442046 470208 442102
rect 469888 441978 470208 442046
rect 469888 441922 469958 441978
rect 470014 441922 470082 441978
rect 470138 441922 470208 441978
rect 469888 441888 470208 441922
rect 500608 442350 500928 442384
rect 500608 442294 500678 442350
rect 500734 442294 500802 442350
rect 500858 442294 500928 442350
rect 500608 442226 500928 442294
rect 500608 442170 500678 442226
rect 500734 442170 500802 442226
rect 500858 442170 500928 442226
rect 500608 442102 500928 442170
rect 500608 442046 500678 442102
rect 500734 442046 500802 442102
rect 500858 442046 500928 442102
rect 500608 441978 500928 442046
rect 500608 441922 500678 441978
rect 500734 441922 500802 441978
rect 500858 441922 500928 441978
rect 500608 441888 500928 441922
rect 24448 436350 24768 436384
rect 24448 436294 24518 436350
rect 24574 436294 24642 436350
rect 24698 436294 24768 436350
rect 24448 436226 24768 436294
rect 24448 436170 24518 436226
rect 24574 436170 24642 436226
rect 24698 436170 24768 436226
rect 24448 436102 24768 436170
rect 24448 436046 24518 436102
rect 24574 436046 24642 436102
rect 24698 436046 24768 436102
rect 24448 435978 24768 436046
rect 24448 435922 24518 435978
rect 24574 435922 24642 435978
rect 24698 435922 24768 435978
rect 24448 435888 24768 435922
rect 55168 436350 55488 436384
rect 55168 436294 55238 436350
rect 55294 436294 55362 436350
rect 55418 436294 55488 436350
rect 55168 436226 55488 436294
rect 55168 436170 55238 436226
rect 55294 436170 55362 436226
rect 55418 436170 55488 436226
rect 55168 436102 55488 436170
rect 55168 436046 55238 436102
rect 55294 436046 55362 436102
rect 55418 436046 55488 436102
rect 55168 435978 55488 436046
rect 55168 435922 55238 435978
rect 55294 435922 55362 435978
rect 55418 435922 55488 435978
rect 55168 435888 55488 435922
rect 85888 436350 86208 436384
rect 85888 436294 85958 436350
rect 86014 436294 86082 436350
rect 86138 436294 86208 436350
rect 85888 436226 86208 436294
rect 85888 436170 85958 436226
rect 86014 436170 86082 436226
rect 86138 436170 86208 436226
rect 85888 436102 86208 436170
rect 85888 436046 85958 436102
rect 86014 436046 86082 436102
rect 86138 436046 86208 436102
rect 85888 435978 86208 436046
rect 85888 435922 85958 435978
rect 86014 435922 86082 435978
rect 86138 435922 86208 435978
rect 85888 435888 86208 435922
rect 116608 436350 116928 436384
rect 116608 436294 116678 436350
rect 116734 436294 116802 436350
rect 116858 436294 116928 436350
rect 116608 436226 116928 436294
rect 116608 436170 116678 436226
rect 116734 436170 116802 436226
rect 116858 436170 116928 436226
rect 116608 436102 116928 436170
rect 116608 436046 116678 436102
rect 116734 436046 116802 436102
rect 116858 436046 116928 436102
rect 116608 435978 116928 436046
rect 116608 435922 116678 435978
rect 116734 435922 116802 435978
rect 116858 435922 116928 435978
rect 116608 435888 116928 435922
rect 147328 436350 147648 436384
rect 147328 436294 147398 436350
rect 147454 436294 147522 436350
rect 147578 436294 147648 436350
rect 147328 436226 147648 436294
rect 147328 436170 147398 436226
rect 147454 436170 147522 436226
rect 147578 436170 147648 436226
rect 147328 436102 147648 436170
rect 147328 436046 147398 436102
rect 147454 436046 147522 436102
rect 147578 436046 147648 436102
rect 147328 435978 147648 436046
rect 147328 435922 147398 435978
rect 147454 435922 147522 435978
rect 147578 435922 147648 435978
rect 147328 435888 147648 435922
rect 178048 436350 178368 436384
rect 178048 436294 178118 436350
rect 178174 436294 178242 436350
rect 178298 436294 178368 436350
rect 178048 436226 178368 436294
rect 178048 436170 178118 436226
rect 178174 436170 178242 436226
rect 178298 436170 178368 436226
rect 178048 436102 178368 436170
rect 178048 436046 178118 436102
rect 178174 436046 178242 436102
rect 178298 436046 178368 436102
rect 178048 435978 178368 436046
rect 178048 435922 178118 435978
rect 178174 435922 178242 435978
rect 178298 435922 178368 435978
rect 178048 435888 178368 435922
rect 208768 436350 209088 436384
rect 208768 436294 208838 436350
rect 208894 436294 208962 436350
rect 209018 436294 209088 436350
rect 208768 436226 209088 436294
rect 208768 436170 208838 436226
rect 208894 436170 208962 436226
rect 209018 436170 209088 436226
rect 208768 436102 209088 436170
rect 208768 436046 208838 436102
rect 208894 436046 208962 436102
rect 209018 436046 209088 436102
rect 208768 435978 209088 436046
rect 208768 435922 208838 435978
rect 208894 435922 208962 435978
rect 209018 435922 209088 435978
rect 208768 435888 209088 435922
rect 239488 436350 239808 436384
rect 239488 436294 239558 436350
rect 239614 436294 239682 436350
rect 239738 436294 239808 436350
rect 239488 436226 239808 436294
rect 239488 436170 239558 436226
rect 239614 436170 239682 436226
rect 239738 436170 239808 436226
rect 239488 436102 239808 436170
rect 239488 436046 239558 436102
rect 239614 436046 239682 436102
rect 239738 436046 239808 436102
rect 239488 435978 239808 436046
rect 239488 435922 239558 435978
rect 239614 435922 239682 435978
rect 239738 435922 239808 435978
rect 239488 435888 239808 435922
rect 270208 436350 270528 436384
rect 270208 436294 270278 436350
rect 270334 436294 270402 436350
rect 270458 436294 270528 436350
rect 270208 436226 270528 436294
rect 270208 436170 270278 436226
rect 270334 436170 270402 436226
rect 270458 436170 270528 436226
rect 270208 436102 270528 436170
rect 270208 436046 270278 436102
rect 270334 436046 270402 436102
rect 270458 436046 270528 436102
rect 270208 435978 270528 436046
rect 270208 435922 270278 435978
rect 270334 435922 270402 435978
rect 270458 435922 270528 435978
rect 270208 435888 270528 435922
rect 300928 436350 301248 436384
rect 300928 436294 300998 436350
rect 301054 436294 301122 436350
rect 301178 436294 301248 436350
rect 300928 436226 301248 436294
rect 300928 436170 300998 436226
rect 301054 436170 301122 436226
rect 301178 436170 301248 436226
rect 300928 436102 301248 436170
rect 300928 436046 300998 436102
rect 301054 436046 301122 436102
rect 301178 436046 301248 436102
rect 300928 435978 301248 436046
rect 300928 435922 300998 435978
rect 301054 435922 301122 435978
rect 301178 435922 301248 435978
rect 300928 435888 301248 435922
rect 331648 436350 331968 436384
rect 331648 436294 331718 436350
rect 331774 436294 331842 436350
rect 331898 436294 331968 436350
rect 331648 436226 331968 436294
rect 331648 436170 331718 436226
rect 331774 436170 331842 436226
rect 331898 436170 331968 436226
rect 331648 436102 331968 436170
rect 331648 436046 331718 436102
rect 331774 436046 331842 436102
rect 331898 436046 331968 436102
rect 331648 435978 331968 436046
rect 331648 435922 331718 435978
rect 331774 435922 331842 435978
rect 331898 435922 331968 435978
rect 331648 435888 331968 435922
rect 362368 436350 362688 436384
rect 362368 436294 362438 436350
rect 362494 436294 362562 436350
rect 362618 436294 362688 436350
rect 362368 436226 362688 436294
rect 362368 436170 362438 436226
rect 362494 436170 362562 436226
rect 362618 436170 362688 436226
rect 362368 436102 362688 436170
rect 362368 436046 362438 436102
rect 362494 436046 362562 436102
rect 362618 436046 362688 436102
rect 362368 435978 362688 436046
rect 362368 435922 362438 435978
rect 362494 435922 362562 435978
rect 362618 435922 362688 435978
rect 362368 435888 362688 435922
rect 393088 436350 393408 436384
rect 393088 436294 393158 436350
rect 393214 436294 393282 436350
rect 393338 436294 393408 436350
rect 393088 436226 393408 436294
rect 393088 436170 393158 436226
rect 393214 436170 393282 436226
rect 393338 436170 393408 436226
rect 393088 436102 393408 436170
rect 393088 436046 393158 436102
rect 393214 436046 393282 436102
rect 393338 436046 393408 436102
rect 393088 435978 393408 436046
rect 393088 435922 393158 435978
rect 393214 435922 393282 435978
rect 393338 435922 393408 435978
rect 393088 435888 393408 435922
rect 423808 436350 424128 436384
rect 423808 436294 423878 436350
rect 423934 436294 424002 436350
rect 424058 436294 424128 436350
rect 423808 436226 424128 436294
rect 423808 436170 423878 436226
rect 423934 436170 424002 436226
rect 424058 436170 424128 436226
rect 423808 436102 424128 436170
rect 423808 436046 423878 436102
rect 423934 436046 424002 436102
rect 424058 436046 424128 436102
rect 423808 435978 424128 436046
rect 423808 435922 423878 435978
rect 423934 435922 424002 435978
rect 424058 435922 424128 435978
rect 423808 435888 424128 435922
rect 454528 436350 454848 436384
rect 454528 436294 454598 436350
rect 454654 436294 454722 436350
rect 454778 436294 454848 436350
rect 454528 436226 454848 436294
rect 454528 436170 454598 436226
rect 454654 436170 454722 436226
rect 454778 436170 454848 436226
rect 454528 436102 454848 436170
rect 454528 436046 454598 436102
rect 454654 436046 454722 436102
rect 454778 436046 454848 436102
rect 454528 435978 454848 436046
rect 454528 435922 454598 435978
rect 454654 435922 454722 435978
rect 454778 435922 454848 435978
rect 454528 435888 454848 435922
rect 485248 436350 485568 436384
rect 485248 436294 485318 436350
rect 485374 436294 485442 436350
rect 485498 436294 485568 436350
rect 485248 436226 485568 436294
rect 485248 436170 485318 436226
rect 485374 436170 485442 436226
rect 485498 436170 485568 436226
rect 485248 436102 485568 436170
rect 485248 436046 485318 436102
rect 485374 436046 485442 436102
rect 485498 436046 485568 436102
rect 485248 435978 485568 436046
rect 485248 435922 485318 435978
rect 485374 435922 485442 435978
rect 485498 435922 485568 435978
rect 485248 435888 485568 435922
rect 515968 436350 516288 436384
rect 515968 436294 516038 436350
rect 516094 436294 516162 436350
rect 516218 436294 516288 436350
rect 515968 436226 516288 436294
rect 515968 436170 516038 436226
rect 516094 436170 516162 436226
rect 516218 436170 516288 436226
rect 515968 436102 516288 436170
rect 515968 436046 516038 436102
rect 516094 436046 516162 436102
rect 516218 436046 516288 436102
rect 515968 435978 516288 436046
rect 515968 435922 516038 435978
rect 516094 435922 516162 435978
rect 516218 435922 516288 435978
rect 515968 435888 516288 435922
rect 525154 436350 525774 453922
rect 525154 436294 525250 436350
rect 525306 436294 525374 436350
rect 525430 436294 525498 436350
rect 525554 436294 525622 436350
rect 525678 436294 525774 436350
rect 525154 436226 525774 436294
rect 525154 436170 525250 436226
rect 525306 436170 525374 436226
rect 525430 436170 525498 436226
rect 525554 436170 525622 436226
rect 525678 436170 525774 436226
rect 525154 436102 525774 436170
rect 525154 436046 525250 436102
rect 525306 436046 525374 436102
rect 525430 436046 525498 436102
rect 525554 436046 525622 436102
rect 525678 436046 525774 436102
rect 525154 435978 525774 436046
rect 525154 435922 525250 435978
rect 525306 435922 525374 435978
rect 525430 435922 525498 435978
rect 525554 435922 525622 435978
rect 525678 435922 525774 435978
rect 6874 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 7494 424350
rect 6874 424226 7494 424294
rect 6874 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 7494 424226
rect 6874 424102 7494 424170
rect 6874 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 7494 424102
rect 6874 423978 7494 424046
rect 6874 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 7494 423978
rect 6874 406350 7494 423922
rect 39808 424350 40128 424384
rect 39808 424294 39878 424350
rect 39934 424294 40002 424350
rect 40058 424294 40128 424350
rect 39808 424226 40128 424294
rect 39808 424170 39878 424226
rect 39934 424170 40002 424226
rect 40058 424170 40128 424226
rect 39808 424102 40128 424170
rect 39808 424046 39878 424102
rect 39934 424046 40002 424102
rect 40058 424046 40128 424102
rect 39808 423978 40128 424046
rect 39808 423922 39878 423978
rect 39934 423922 40002 423978
rect 40058 423922 40128 423978
rect 39808 423888 40128 423922
rect 70528 424350 70848 424384
rect 70528 424294 70598 424350
rect 70654 424294 70722 424350
rect 70778 424294 70848 424350
rect 70528 424226 70848 424294
rect 70528 424170 70598 424226
rect 70654 424170 70722 424226
rect 70778 424170 70848 424226
rect 70528 424102 70848 424170
rect 70528 424046 70598 424102
rect 70654 424046 70722 424102
rect 70778 424046 70848 424102
rect 70528 423978 70848 424046
rect 70528 423922 70598 423978
rect 70654 423922 70722 423978
rect 70778 423922 70848 423978
rect 70528 423888 70848 423922
rect 101248 424350 101568 424384
rect 101248 424294 101318 424350
rect 101374 424294 101442 424350
rect 101498 424294 101568 424350
rect 101248 424226 101568 424294
rect 101248 424170 101318 424226
rect 101374 424170 101442 424226
rect 101498 424170 101568 424226
rect 101248 424102 101568 424170
rect 101248 424046 101318 424102
rect 101374 424046 101442 424102
rect 101498 424046 101568 424102
rect 101248 423978 101568 424046
rect 101248 423922 101318 423978
rect 101374 423922 101442 423978
rect 101498 423922 101568 423978
rect 101248 423888 101568 423922
rect 131968 424350 132288 424384
rect 131968 424294 132038 424350
rect 132094 424294 132162 424350
rect 132218 424294 132288 424350
rect 131968 424226 132288 424294
rect 131968 424170 132038 424226
rect 132094 424170 132162 424226
rect 132218 424170 132288 424226
rect 131968 424102 132288 424170
rect 131968 424046 132038 424102
rect 132094 424046 132162 424102
rect 132218 424046 132288 424102
rect 131968 423978 132288 424046
rect 131968 423922 132038 423978
rect 132094 423922 132162 423978
rect 132218 423922 132288 423978
rect 131968 423888 132288 423922
rect 162688 424350 163008 424384
rect 162688 424294 162758 424350
rect 162814 424294 162882 424350
rect 162938 424294 163008 424350
rect 162688 424226 163008 424294
rect 162688 424170 162758 424226
rect 162814 424170 162882 424226
rect 162938 424170 163008 424226
rect 162688 424102 163008 424170
rect 162688 424046 162758 424102
rect 162814 424046 162882 424102
rect 162938 424046 163008 424102
rect 162688 423978 163008 424046
rect 162688 423922 162758 423978
rect 162814 423922 162882 423978
rect 162938 423922 163008 423978
rect 162688 423888 163008 423922
rect 193408 424350 193728 424384
rect 193408 424294 193478 424350
rect 193534 424294 193602 424350
rect 193658 424294 193728 424350
rect 193408 424226 193728 424294
rect 193408 424170 193478 424226
rect 193534 424170 193602 424226
rect 193658 424170 193728 424226
rect 193408 424102 193728 424170
rect 193408 424046 193478 424102
rect 193534 424046 193602 424102
rect 193658 424046 193728 424102
rect 193408 423978 193728 424046
rect 193408 423922 193478 423978
rect 193534 423922 193602 423978
rect 193658 423922 193728 423978
rect 193408 423888 193728 423922
rect 224128 424350 224448 424384
rect 224128 424294 224198 424350
rect 224254 424294 224322 424350
rect 224378 424294 224448 424350
rect 224128 424226 224448 424294
rect 224128 424170 224198 424226
rect 224254 424170 224322 424226
rect 224378 424170 224448 424226
rect 224128 424102 224448 424170
rect 224128 424046 224198 424102
rect 224254 424046 224322 424102
rect 224378 424046 224448 424102
rect 224128 423978 224448 424046
rect 224128 423922 224198 423978
rect 224254 423922 224322 423978
rect 224378 423922 224448 423978
rect 224128 423888 224448 423922
rect 254848 424350 255168 424384
rect 254848 424294 254918 424350
rect 254974 424294 255042 424350
rect 255098 424294 255168 424350
rect 254848 424226 255168 424294
rect 254848 424170 254918 424226
rect 254974 424170 255042 424226
rect 255098 424170 255168 424226
rect 254848 424102 255168 424170
rect 254848 424046 254918 424102
rect 254974 424046 255042 424102
rect 255098 424046 255168 424102
rect 254848 423978 255168 424046
rect 254848 423922 254918 423978
rect 254974 423922 255042 423978
rect 255098 423922 255168 423978
rect 254848 423888 255168 423922
rect 285568 424350 285888 424384
rect 285568 424294 285638 424350
rect 285694 424294 285762 424350
rect 285818 424294 285888 424350
rect 285568 424226 285888 424294
rect 285568 424170 285638 424226
rect 285694 424170 285762 424226
rect 285818 424170 285888 424226
rect 285568 424102 285888 424170
rect 285568 424046 285638 424102
rect 285694 424046 285762 424102
rect 285818 424046 285888 424102
rect 285568 423978 285888 424046
rect 285568 423922 285638 423978
rect 285694 423922 285762 423978
rect 285818 423922 285888 423978
rect 285568 423888 285888 423922
rect 316288 424350 316608 424384
rect 316288 424294 316358 424350
rect 316414 424294 316482 424350
rect 316538 424294 316608 424350
rect 316288 424226 316608 424294
rect 316288 424170 316358 424226
rect 316414 424170 316482 424226
rect 316538 424170 316608 424226
rect 316288 424102 316608 424170
rect 316288 424046 316358 424102
rect 316414 424046 316482 424102
rect 316538 424046 316608 424102
rect 316288 423978 316608 424046
rect 316288 423922 316358 423978
rect 316414 423922 316482 423978
rect 316538 423922 316608 423978
rect 316288 423888 316608 423922
rect 347008 424350 347328 424384
rect 347008 424294 347078 424350
rect 347134 424294 347202 424350
rect 347258 424294 347328 424350
rect 347008 424226 347328 424294
rect 347008 424170 347078 424226
rect 347134 424170 347202 424226
rect 347258 424170 347328 424226
rect 347008 424102 347328 424170
rect 347008 424046 347078 424102
rect 347134 424046 347202 424102
rect 347258 424046 347328 424102
rect 347008 423978 347328 424046
rect 347008 423922 347078 423978
rect 347134 423922 347202 423978
rect 347258 423922 347328 423978
rect 347008 423888 347328 423922
rect 377728 424350 378048 424384
rect 377728 424294 377798 424350
rect 377854 424294 377922 424350
rect 377978 424294 378048 424350
rect 377728 424226 378048 424294
rect 377728 424170 377798 424226
rect 377854 424170 377922 424226
rect 377978 424170 378048 424226
rect 377728 424102 378048 424170
rect 377728 424046 377798 424102
rect 377854 424046 377922 424102
rect 377978 424046 378048 424102
rect 377728 423978 378048 424046
rect 377728 423922 377798 423978
rect 377854 423922 377922 423978
rect 377978 423922 378048 423978
rect 377728 423888 378048 423922
rect 408448 424350 408768 424384
rect 408448 424294 408518 424350
rect 408574 424294 408642 424350
rect 408698 424294 408768 424350
rect 408448 424226 408768 424294
rect 408448 424170 408518 424226
rect 408574 424170 408642 424226
rect 408698 424170 408768 424226
rect 408448 424102 408768 424170
rect 408448 424046 408518 424102
rect 408574 424046 408642 424102
rect 408698 424046 408768 424102
rect 408448 423978 408768 424046
rect 408448 423922 408518 423978
rect 408574 423922 408642 423978
rect 408698 423922 408768 423978
rect 408448 423888 408768 423922
rect 439168 424350 439488 424384
rect 439168 424294 439238 424350
rect 439294 424294 439362 424350
rect 439418 424294 439488 424350
rect 439168 424226 439488 424294
rect 439168 424170 439238 424226
rect 439294 424170 439362 424226
rect 439418 424170 439488 424226
rect 439168 424102 439488 424170
rect 439168 424046 439238 424102
rect 439294 424046 439362 424102
rect 439418 424046 439488 424102
rect 439168 423978 439488 424046
rect 439168 423922 439238 423978
rect 439294 423922 439362 423978
rect 439418 423922 439488 423978
rect 439168 423888 439488 423922
rect 469888 424350 470208 424384
rect 469888 424294 469958 424350
rect 470014 424294 470082 424350
rect 470138 424294 470208 424350
rect 469888 424226 470208 424294
rect 469888 424170 469958 424226
rect 470014 424170 470082 424226
rect 470138 424170 470208 424226
rect 469888 424102 470208 424170
rect 469888 424046 469958 424102
rect 470014 424046 470082 424102
rect 470138 424046 470208 424102
rect 469888 423978 470208 424046
rect 469888 423922 469958 423978
rect 470014 423922 470082 423978
rect 470138 423922 470208 423978
rect 469888 423888 470208 423922
rect 500608 424350 500928 424384
rect 500608 424294 500678 424350
rect 500734 424294 500802 424350
rect 500858 424294 500928 424350
rect 500608 424226 500928 424294
rect 500608 424170 500678 424226
rect 500734 424170 500802 424226
rect 500858 424170 500928 424226
rect 500608 424102 500928 424170
rect 500608 424046 500678 424102
rect 500734 424046 500802 424102
rect 500858 424046 500928 424102
rect 500608 423978 500928 424046
rect 500608 423922 500678 423978
rect 500734 423922 500802 423978
rect 500858 423922 500928 423978
rect 500608 423888 500928 423922
rect 24448 418350 24768 418384
rect 24448 418294 24518 418350
rect 24574 418294 24642 418350
rect 24698 418294 24768 418350
rect 24448 418226 24768 418294
rect 24448 418170 24518 418226
rect 24574 418170 24642 418226
rect 24698 418170 24768 418226
rect 24448 418102 24768 418170
rect 24448 418046 24518 418102
rect 24574 418046 24642 418102
rect 24698 418046 24768 418102
rect 24448 417978 24768 418046
rect 24448 417922 24518 417978
rect 24574 417922 24642 417978
rect 24698 417922 24768 417978
rect 24448 417888 24768 417922
rect 55168 418350 55488 418384
rect 55168 418294 55238 418350
rect 55294 418294 55362 418350
rect 55418 418294 55488 418350
rect 55168 418226 55488 418294
rect 55168 418170 55238 418226
rect 55294 418170 55362 418226
rect 55418 418170 55488 418226
rect 55168 418102 55488 418170
rect 55168 418046 55238 418102
rect 55294 418046 55362 418102
rect 55418 418046 55488 418102
rect 55168 417978 55488 418046
rect 55168 417922 55238 417978
rect 55294 417922 55362 417978
rect 55418 417922 55488 417978
rect 55168 417888 55488 417922
rect 85888 418350 86208 418384
rect 85888 418294 85958 418350
rect 86014 418294 86082 418350
rect 86138 418294 86208 418350
rect 85888 418226 86208 418294
rect 85888 418170 85958 418226
rect 86014 418170 86082 418226
rect 86138 418170 86208 418226
rect 85888 418102 86208 418170
rect 85888 418046 85958 418102
rect 86014 418046 86082 418102
rect 86138 418046 86208 418102
rect 85888 417978 86208 418046
rect 85888 417922 85958 417978
rect 86014 417922 86082 417978
rect 86138 417922 86208 417978
rect 85888 417888 86208 417922
rect 116608 418350 116928 418384
rect 116608 418294 116678 418350
rect 116734 418294 116802 418350
rect 116858 418294 116928 418350
rect 116608 418226 116928 418294
rect 116608 418170 116678 418226
rect 116734 418170 116802 418226
rect 116858 418170 116928 418226
rect 116608 418102 116928 418170
rect 116608 418046 116678 418102
rect 116734 418046 116802 418102
rect 116858 418046 116928 418102
rect 116608 417978 116928 418046
rect 116608 417922 116678 417978
rect 116734 417922 116802 417978
rect 116858 417922 116928 417978
rect 116608 417888 116928 417922
rect 147328 418350 147648 418384
rect 147328 418294 147398 418350
rect 147454 418294 147522 418350
rect 147578 418294 147648 418350
rect 147328 418226 147648 418294
rect 147328 418170 147398 418226
rect 147454 418170 147522 418226
rect 147578 418170 147648 418226
rect 147328 418102 147648 418170
rect 147328 418046 147398 418102
rect 147454 418046 147522 418102
rect 147578 418046 147648 418102
rect 147328 417978 147648 418046
rect 147328 417922 147398 417978
rect 147454 417922 147522 417978
rect 147578 417922 147648 417978
rect 147328 417888 147648 417922
rect 178048 418350 178368 418384
rect 178048 418294 178118 418350
rect 178174 418294 178242 418350
rect 178298 418294 178368 418350
rect 178048 418226 178368 418294
rect 178048 418170 178118 418226
rect 178174 418170 178242 418226
rect 178298 418170 178368 418226
rect 178048 418102 178368 418170
rect 178048 418046 178118 418102
rect 178174 418046 178242 418102
rect 178298 418046 178368 418102
rect 178048 417978 178368 418046
rect 178048 417922 178118 417978
rect 178174 417922 178242 417978
rect 178298 417922 178368 417978
rect 178048 417888 178368 417922
rect 208768 418350 209088 418384
rect 208768 418294 208838 418350
rect 208894 418294 208962 418350
rect 209018 418294 209088 418350
rect 208768 418226 209088 418294
rect 208768 418170 208838 418226
rect 208894 418170 208962 418226
rect 209018 418170 209088 418226
rect 208768 418102 209088 418170
rect 208768 418046 208838 418102
rect 208894 418046 208962 418102
rect 209018 418046 209088 418102
rect 208768 417978 209088 418046
rect 208768 417922 208838 417978
rect 208894 417922 208962 417978
rect 209018 417922 209088 417978
rect 208768 417888 209088 417922
rect 239488 418350 239808 418384
rect 239488 418294 239558 418350
rect 239614 418294 239682 418350
rect 239738 418294 239808 418350
rect 239488 418226 239808 418294
rect 239488 418170 239558 418226
rect 239614 418170 239682 418226
rect 239738 418170 239808 418226
rect 239488 418102 239808 418170
rect 239488 418046 239558 418102
rect 239614 418046 239682 418102
rect 239738 418046 239808 418102
rect 239488 417978 239808 418046
rect 239488 417922 239558 417978
rect 239614 417922 239682 417978
rect 239738 417922 239808 417978
rect 239488 417888 239808 417922
rect 270208 418350 270528 418384
rect 270208 418294 270278 418350
rect 270334 418294 270402 418350
rect 270458 418294 270528 418350
rect 270208 418226 270528 418294
rect 270208 418170 270278 418226
rect 270334 418170 270402 418226
rect 270458 418170 270528 418226
rect 270208 418102 270528 418170
rect 270208 418046 270278 418102
rect 270334 418046 270402 418102
rect 270458 418046 270528 418102
rect 270208 417978 270528 418046
rect 270208 417922 270278 417978
rect 270334 417922 270402 417978
rect 270458 417922 270528 417978
rect 270208 417888 270528 417922
rect 300928 418350 301248 418384
rect 300928 418294 300998 418350
rect 301054 418294 301122 418350
rect 301178 418294 301248 418350
rect 300928 418226 301248 418294
rect 300928 418170 300998 418226
rect 301054 418170 301122 418226
rect 301178 418170 301248 418226
rect 300928 418102 301248 418170
rect 300928 418046 300998 418102
rect 301054 418046 301122 418102
rect 301178 418046 301248 418102
rect 300928 417978 301248 418046
rect 300928 417922 300998 417978
rect 301054 417922 301122 417978
rect 301178 417922 301248 417978
rect 300928 417888 301248 417922
rect 331648 418350 331968 418384
rect 331648 418294 331718 418350
rect 331774 418294 331842 418350
rect 331898 418294 331968 418350
rect 331648 418226 331968 418294
rect 331648 418170 331718 418226
rect 331774 418170 331842 418226
rect 331898 418170 331968 418226
rect 331648 418102 331968 418170
rect 331648 418046 331718 418102
rect 331774 418046 331842 418102
rect 331898 418046 331968 418102
rect 331648 417978 331968 418046
rect 331648 417922 331718 417978
rect 331774 417922 331842 417978
rect 331898 417922 331968 417978
rect 331648 417888 331968 417922
rect 362368 418350 362688 418384
rect 362368 418294 362438 418350
rect 362494 418294 362562 418350
rect 362618 418294 362688 418350
rect 362368 418226 362688 418294
rect 362368 418170 362438 418226
rect 362494 418170 362562 418226
rect 362618 418170 362688 418226
rect 362368 418102 362688 418170
rect 362368 418046 362438 418102
rect 362494 418046 362562 418102
rect 362618 418046 362688 418102
rect 362368 417978 362688 418046
rect 362368 417922 362438 417978
rect 362494 417922 362562 417978
rect 362618 417922 362688 417978
rect 362368 417888 362688 417922
rect 393088 418350 393408 418384
rect 393088 418294 393158 418350
rect 393214 418294 393282 418350
rect 393338 418294 393408 418350
rect 393088 418226 393408 418294
rect 393088 418170 393158 418226
rect 393214 418170 393282 418226
rect 393338 418170 393408 418226
rect 393088 418102 393408 418170
rect 393088 418046 393158 418102
rect 393214 418046 393282 418102
rect 393338 418046 393408 418102
rect 393088 417978 393408 418046
rect 393088 417922 393158 417978
rect 393214 417922 393282 417978
rect 393338 417922 393408 417978
rect 393088 417888 393408 417922
rect 423808 418350 424128 418384
rect 423808 418294 423878 418350
rect 423934 418294 424002 418350
rect 424058 418294 424128 418350
rect 423808 418226 424128 418294
rect 423808 418170 423878 418226
rect 423934 418170 424002 418226
rect 424058 418170 424128 418226
rect 423808 418102 424128 418170
rect 423808 418046 423878 418102
rect 423934 418046 424002 418102
rect 424058 418046 424128 418102
rect 423808 417978 424128 418046
rect 423808 417922 423878 417978
rect 423934 417922 424002 417978
rect 424058 417922 424128 417978
rect 423808 417888 424128 417922
rect 454528 418350 454848 418384
rect 454528 418294 454598 418350
rect 454654 418294 454722 418350
rect 454778 418294 454848 418350
rect 454528 418226 454848 418294
rect 454528 418170 454598 418226
rect 454654 418170 454722 418226
rect 454778 418170 454848 418226
rect 454528 418102 454848 418170
rect 454528 418046 454598 418102
rect 454654 418046 454722 418102
rect 454778 418046 454848 418102
rect 454528 417978 454848 418046
rect 454528 417922 454598 417978
rect 454654 417922 454722 417978
rect 454778 417922 454848 417978
rect 454528 417888 454848 417922
rect 485248 418350 485568 418384
rect 485248 418294 485318 418350
rect 485374 418294 485442 418350
rect 485498 418294 485568 418350
rect 485248 418226 485568 418294
rect 485248 418170 485318 418226
rect 485374 418170 485442 418226
rect 485498 418170 485568 418226
rect 485248 418102 485568 418170
rect 485248 418046 485318 418102
rect 485374 418046 485442 418102
rect 485498 418046 485568 418102
rect 485248 417978 485568 418046
rect 485248 417922 485318 417978
rect 485374 417922 485442 417978
rect 485498 417922 485568 417978
rect 485248 417888 485568 417922
rect 515968 418350 516288 418384
rect 515968 418294 516038 418350
rect 516094 418294 516162 418350
rect 516218 418294 516288 418350
rect 515968 418226 516288 418294
rect 515968 418170 516038 418226
rect 516094 418170 516162 418226
rect 516218 418170 516288 418226
rect 515968 418102 516288 418170
rect 515968 418046 516038 418102
rect 516094 418046 516162 418102
rect 516218 418046 516288 418102
rect 515968 417978 516288 418046
rect 515968 417922 516038 417978
rect 516094 417922 516162 417978
rect 516218 417922 516288 417978
rect 515968 417888 516288 417922
rect 525154 418350 525774 435922
rect 525154 418294 525250 418350
rect 525306 418294 525374 418350
rect 525430 418294 525498 418350
rect 525554 418294 525622 418350
rect 525678 418294 525774 418350
rect 525154 418226 525774 418294
rect 525154 418170 525250 418226
rect 525306 418170 525374 418226
rect 525430 418170 525498 418226
rect 525554 418170 525622 418226
rect 525678 418170 525774 418226
rect 525154 418102 525774 418170
rect 525154 418046 525250 418102
rect 525306 418046 525374 418102
rect 525430 418046 525498 418102
rect 525554 418046 525622 418102
rect 525678 418046 525774 418102
rect 525154 417978 525774 418046
rect 525154 417922 525250 417978
rect 525306 417922 525374 417978
rect 525430 417922 525498 417978
rect 525554 417922 525622 417978
rect 525678 417922 525774 417978
rect 6874 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 7494 406350
rect 6874 406226 7494 406294
rect 6874 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 7494 406226
rect 6874 406102 7494 406170
rect 6874 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 7494 406102
rect 6874 405978 7494 406046
rect 6874 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 7494 405978
rect 6874 388350 7494 405922
rect 39808 406350 40128 406384
rect 39808 406294 39878 406350
rect 39934 406294 40002 406350
rect 40058 406294 40128 406350
rect 39808 406226 40128 406294
rect 39808 406170 39878 406226
rect 39934 406170 40002 406226
rect 40058 406170 40128 406226
rect 39808 406102 40128 406170
rect 39808 406046 39878 406102
rect 39934 406046 40002 406102
rect 40058 406046 40128 406102
rect 39808 405978 40128 406046
rect 39808 405922 39878 405978
rect 39934 405922 40002 405978
rect 40058 405922 40128 405978
rect 39808 405888 40128 405922
rect 70528 406350 70848 406384
rect 70528 406294 70598 406350
rect 70654 406294 70722 406350
rect 70778 406294 70848 406350
rect 70528 406226 70848 406294
rect 70528 406170 70598 406226
rect 70654 406170 70722 406226
rect 70778 406170 70848 406226
rect 70528 406102 70848 406170
rect 70528 406046 70598 406102
rect 70654 406046 70722 406102
rect 70778 406046 70848 406102
rect 70528 405978 70848 406046
rect 70528 405922 70598 405978
rect 70654 405922 70722 405978
rect 70778 405922 70848 405978
rect 70528 405888 70848 405922
rect 101248 406350 101568 406384
rect 101248 406294 101318 406350
rect 101374 406294 101442 406350
rect 101498 406294 101568 406350
rect 101248 406226 101568 406294
rect 101248 406170 101318 406226
rect 101374 406170 101442 406226
rect 101498 406170 101568 406226
rect 101248 406102 101568 406170
rect 101248 406046 101318 406102
rect 101374 406046 101442 406102
rect 101498 406046 101568 406102
rect 101248 405978 101568 406046
rect 101248 405922 101318 405978
rect 101374 405922 101442 405978
rect 101498 405922 101568 405978
rect 101248 405888 101568 405922
rect 131968 406350 132288 406384
rect 131968 406294 132038 406350
rect 132094 406294 132162 406350
rect 132218 406294 132288 406350
rect 131968 406226 132288 406294
rect 131968 406170 132038 406226
rect 132094 406170 132162 406226
rect 132218 406170 132288 406226
rect 131968 406102 132288 406170
rect 131968 406046 132038 406102
rect 132094 406046 132162 406102
rect 132218 406046 132288 406102
rect 131968 405978 132288 406046
rect 131968 405922 132038 405978
rect 132094 405922 132162 405978
rect 132218 405922 132288 405978
rect 131968 405888 132288 405922
rect 162688 406350 163008 406384
rect 162688 406294 162758 406350
rect 162814 406294 162882 406350
rect 162938 406294 163008 406350
rect 162688 406226 163008 406294
rect 162688 406170 162758 406226
rect 162814 406170 162882 406226
rect 162938 406170 163008 406226
rect 162688 406102 163008 406170
rect 162688 406046 162758 406102
rect 162814 406046 162882 406102
rect 162938 406046 163008 406102
rect 162688 405978 163008 406046
rect 162688 405922 162758 405978
rect 162814 405922 162882 405978
rect 162938 405922 163008 405978
rect 162688 405888 163008 405922
rect 193408 406350 193728 406384
rect 193408 406294 193478 406350
rect 193534 406294 193602 406350
rect 193658 406294 193728 406350
rect 193408 406226 193728 406294
rect 193408 406170 193478 406226
rect 193534 406170 193602 406226
rect 193658 406170 193728 406226
rect 193408 406102 193728 406170
rect 193408 406046 193478 406102
rect 193534 406046 193602 406102
rect 193658 406046 193728 406102
rect 193408 405978 193728 406046
rect 193408 405922 193478 405978
rect 193534 405922 193602 405978
rect 193658 405922 193728 405978
rect 193408 405888 193728 405922
rect 224128 406350 224448 406384
rect 224128 406294 224198 406350
rect 224254 406294 224322 406350
rect 224378 406294 224448 406350
rect 224128 406226 224448 406294
rect 224128 406170 224198 406226
rect 224254 406170 224322 406226
rect 224378 406170 224448 406226
rect 224128 406102 224448 406170
rect 224128 406046 224198 406102
rect 224254 406046 224322 406102
rect 224378 406046 224448 406102
rect 224128 405978 224448 406046
rect 224128 405922 224198 405978
rect 224254 405922 224322 405978
rect 224378 405922 224448 405978
rect 224128 405888 224448 405922
rect 254848 406350 255168 406384
rect 254848 406294 254918 406350
rect 254974 406294 255042 406350
rect 255098 406294 255168 406350
rect 254848 406226 255168 406294
rect 254848 406170 254918 406226
rect 254974 406170 255042 406226
rect 255098 406170 255168 406226
rect 254848 406102 255168 406170
rect 254848 406046 254918 406102
rect 254974 406046 255042 406102
rect 255098 406046 255168 406102
rect 254848 405978 255168 406046
rect 254848 405922 254918 405978
rect 254974 405922 255042 405978
rect 255098 405922 255168 405978
rect 254848 405888 255168 405922
rect 285568 406350 285888 406384
rect 285568 406294 285638 406350
rect 285694 406294 285762 406350
rect 285818 406294 285888 406350
rect 285568 406226 285888 406294
rect 285568 406170 285638 406226
rect 285694 406170 285762 406226
rect 285818 406170 285888 406226
rect 285568 406102 285888 406170
rect 285568 406046 285638 406102
rect 285694 406046 285762 406102
rect 285818 406046 285888 406102
rect 285568 405978 285888 406046
rect 285568 405922 285638 405978
rect 285694 405922 285762 405978
rect 285818 405922 285888 405978
rect 285568 405888 285888 405922
rect 316288 406350 316608 406384
rect 316288 406294 316358 406350
rect 316414 406294 316482 406350
rect 316538 406294 316608 406350
rect 316288 406226 316608 406294
rect 316288 406170 316358 406226
rect 316414 406170 316482 406226
rect 316538 406170 316608 406226
rect 316288 406102 316608 406170
rect 316288 406046 316358 406102
rect 316414 406046 316482 406102
rect 316538 406046 316608 406102
rect 316288 405978 316608 406046
rect 316288 405922 316358 405978
rect 316414 405922 316482 405978
rect 316538 405922 316608 405978
rect 316288 405888 316608 405922
rect 347008 406350 347328 406384
rect 347008 406294 347078 406350
rect 347134 406294 347202 406350
rect 347258 406294 347328 406350
rect 347008 406226 347328 406294
rect 347008 406170 347078 406226
rect 347134 406170 347202 406226
rect 347258 406170 347328 406226
rect 347008 406102 347328 406170
rect 347008 406046 347078 406102
rect 347134 406046 347202 406102
rect 347258 406046 347328 406102
rect 347008 405978 347328 406046
rect 347008 405922 347078 405978
rect 347134 405922 347202 405978
rect 347258 405922 347328 405978
rect 347008 405888 347328 405922
rect 377728 406350 378048 406384
rect 377728 406294 377798 406350
rect 377854 406294 377922 406350
rect 377978 406294 378048 406350
rect 377728 406226 378048 406294
rect 377728 406170 377798 406226
rect 377854 406170 377922 406226
rect 377978 406170 378048 406226
rect 377728 406102 378048 406170
rect 377728 406046 377798 406102
rect 377854 406046 377922 406102
rect 377978 406046 378048 406102
rect 377728 405978 378048 406046
rect 377728 405922 377798 405978
rect 377854 405922 377922 405978
rect 377978 405922 378048 405978
rect 377728 405888 378048 405922
rect 408448 406350 408768 406384
rect 408448 406294 408518 406350
rect 408574 406294 408642 406350
rect 408698 406294 408768 406350
rect 408448 406226 408768 406294
rect 408448 406170 408518 406226
rect 408574 406170 408642 406226
rect 408698 406170 408768 406226
rect 408448 406102 408768 406170
rect 408448 406046 408518 406102
rect 408574 406046 408642 406102
rect 408698 406046 408768 406102
rect 408448 405978 408768 406046
rect 408448 405922 408518 405978
rect 408574 405922 408642 405978
rect 408698 405922 408768 405978
rect 408448 405888 408768 405922
rect 439168 406350 439488 406384
rect 439168 406294 439238 406350
rect 439294 406294 439362 406350
rect 439418 406294 439488 406350
rect 439168 406226 439488 406294
rect 439168 406170 439238 406226
rect 439294 406170 439362 406226
rect 439418 406170 439488 406226
rect 439168 406102 439488 406170
rect 439168 406046 439238 406102
rect 439294 406046 439362 406102
rect 439418 406046 439488 406102
rect 439168 405978 439488 406046
rect 439168 405922 439238 405978
rect 439294 405922 439362 405978
rect 439418 405922 439488 405978
rect 439168 405888 439488 405922
rect 469888 406350 470208 406384
rect 469888 406294 469958 406350
rect 470014 406294 470082 406350
rect 470138 406294 470208 406350
rect 469888 406226 470208 406294
rect 469888 406170 469958 406226
rect 470014 406170 470082 406226
rect 470138 406170 470208 406226
rect 469888 406102 470208 406170
rect 469888 406046 469958 406102
rect 470014 406046 470082 406102
rect 470138 406046 470208 406102
rect 469888 405978 470208 406046
rect 469888 405922 469958 405978
rect 470014 405922 470082 405978
rect 470138 405922 470208 405978
rect 469888 405888 470208 405922
rect 500608 406350 500928 406384
rect 500608 406294 500678 406350
rect 500734 406294 500802 406350
rect 500858 406294 500928 406350
rect 500608 406226 500928 406294
rect 500608 406170 500678 406226
rect 500734 406170 500802 406226
rect 500858 406170 500928 406226
rect 500608 406102 500928 406170
rect 500608 406046 500678 406102
rect 500734 406046 500802 406102
rect 500858 406046 500928 406102
rect 500608 405978 500928 406046
rect 500608 405922 500678 405978
rect 500734 405922 500802 405978
rect 500858 405922 500928 405978
rect 500608 405888 500928 405922
rect 24448 400350 24768 400384
rect 24448 400294 24518 400350
rect 24574 400294 24642 400350
rect 24698 400294 24768 400350
rect 24448 400226 24768 400294
rect 24448 400170 24518 400226
rect 24574 400170 24642 400226
rect 24698 400170 24768 400226
rect 24448 400102 24768 400170
rect 24448 400046 24518 400102
rect 24574 400046 24642 400102
rect 24698 400046 24768 400102
rect 24448 399978 24768 400046
rect 24448 399922 24518 399978
rect 24574 399922 24642 399978
rect 24698 399922 24768 399978
rect 24448 399888 24768 399922
rect 55168 400350 55488 400384
rect 55168 400294 55238 400350
rect 55294 400294 55362 400350
rect 55418 400294 55488 400350
rect 55168 400226 55488 400294
rect 55168 400170 55238 400226
rect 55294 400170 55362 400226
rect 55418 400170 55488 400226
rect 55168 400102 55488 400170
rect 55168 400046 55238 400102
rect 55294 400046 55362 400102
rect 55418 400046 55488 400102
rect 55168 399978 55488 400046
rect 55168 399922 55238 399978
rect 55294 399922 55362 399978
rect 55418 399922 55488 399978
rect 55168 399888 55488 399922
rect 85888 400350 86208 400384
rect 85888 400294 85958 400350
rect 86014 400294 86082 400350
rect 86138 400294 86208 400350
rect 85888 400226 86208 400294
rect 85888 400170 85958 400226
rect 86014 400170 86082 400226
rect 86138 400170 86208 400226
rect 85888 400102 86208 400170
rect 85888 400046 85958 400102
rect 86014 400046 86082 400102
rect 86138 400046 86208 400102
rect 85888 399978 86208 400046
rect 85888 399922 85958 399978
rect 86014 399922 86082 399978
rect 86138 399922 86208 399978
rect 85888 399888 86208 399922
rect 116608 400350 116928 400384
rect 116608 400294 116678 400350
rect 116734 400294 116802 400350
rect 116858 400294 116928 400350
rect 116608 400226 116928 400294
rect 116608 400170 116678 400226
rect 116734 400170 116802 400226
rect 116858 400170 116928 400226
rect 116608 400102 116928 400170
rect 116608 400046 116678 400102
rect 116734 400046 116802 400102
rect 116858 400046 116928 400102
rect 116608 399978 116928 400046
rect 116608 399922 116678 399978
rect 116734 399922 116802 399978
rect 116858 399922 116928 399978
rect 116608 399888 116928 399922
rect 147328 400350 147648 400384
rect 147328 400294 147398 400350
rect 147454 400294 147522 400350
rect 147578 400294 147648 400350
rect 147328 400226 147648 400294
rect 147328 400170 147398 400226
rect 147454 400170 147522 400226
rect 147578 400170 147648 400226
rect 147328 400102 147648 400170
rect 147328 400046 147398 400102
rect 147454 400046 147522 400102
rect 147578 400046 147648 400102
rect 147328 399978 147648 400046
rect 147328 399922 147398 399978
rect 147454 399922 147522 399978
rect 147578 399922 147648 399978
rect 147328 399888 147648 399922
rect 178048 400350 178368 400384
rect 178048 400294 178118 400350
rect 178174 400294 178242 400350
rect 178298 400294 178368 400350
rect 178048 400226 178368 400294
rect 178048 400170 178118 400226
rect 178174 400170 178242 400226
rect 178298 400170 178368 400226
rect 178048 400102 178368 400170
rect 178048 400046 178118 400102
rect 178174 400046 178242 400102
rect 178298 400046 178368 400102
rect 178048 399978 178368 400046
rect 178048 399922 178118 399978
rect 178174 399922 178242 399978
rect 178298 399922 178368 399978
rect 178048 399888 178368 399922
rect 208768 400350 209088 400384
rect 208768 400294 208838 400350
rect 208894 400294 208962 400350
rect 209018 400294 209088 400350
rect 208768 400226 209088 400294
rect 208768 400170 208838 400226
rect 208894 400170 208962 400226
rect 209018 400170 209088 400226
rect 208768 400102 209088 400170
rect 208768 400046 208838 400102
rect 208894 400046 208962 400102
rect 209018 400046 209088 400102
rect 208768 399978 209088 400046
rect 208768 399922 208838 399978
rect 208894 399922 208962 399978
rect 209018 399922 209088 399978
rect 208768 399888 209088 399922
rect 239488 400350 239808 400384
rect 239488 400294 239558 400350
rect 239614 400294 239682 400350
rect 239738 400294 239808 400350
rect 239488 400226 239808 400294
rect 239488 400170 239558 400226
rect 239614 400170 239682 400226
rect 239738 400170 239808 400226
rect 239488 400102 239808 400170
rect 239488 400046 239558 400102
rect 239614 400046 239682 400102
rect 239738 400046 239808 400102
rect 239488 399978 239808 400046
rect 239488 399922 239558 399978
rect 239614 399922 239682 399978
rect 239738 399922 239808 399978
rect 239488 399888 239808 399922
rect 270208 400350 270528 400384
rect 270208 400294 270278 400350
rect 270334 400294 270402 400350
rect 270458 400294 270528 400350
rect 270208 400226 270528 400294
rect 270208 400170 270278 400226
rect 270334 400170 270402 400226
rect 270458 400170 270528 400226
rect 270208 400102 270528 400170
rect 270208 400046 270278 400102
rect 270334 400046 270402 400102
rect 270458 400046 270528 400102
rect 270208 399978 270528 400046
rect 270208 399922 270278 399978
rect 270334 399922 270402 399978
rect 270458 399922 270528 399978
rect 270208 399888 270528 399922
rect 300928 400350 301248 400384
rect 300928 400294 300998 400350
rect 301054 400294 301122 400350
rect 301178 400294 301248 400350
rect 300928 400226 301248 400294
rect 300928 400170 300998 400226
rect 301054 400170 301122 400226
rect 301178 400170 301248 400226
rect 300928 400102 301248 400170
rect 300928 400046 300998 400102
rect 301054 400046 301122 400102
rect 301178 400046 301248 400102
rect 300928 399978 301248 400046
rect 300928 399922 300998 399978
rect 301054 399922 301122 399978
rect 301178 399922 301248 399978
rect 300928 399888 301248 399922
rect 331648 400350 331968 400384
rect 331648 400294 331718 400350
rect 331774 400294 331842 400350
rect 331898 400294 331968 400350
rect 331648 400226 331968 400294
rect 331648 400170 331718 400226
rect 331774 400170 331842 400226
rect 331898 400170 331968 400226
rect 331648 400102 331968 400170
rect 331648 400046 331718 400102
rect 331774 400046 331842 400102
rect 331898 400046 331968 400102
rect 331648 399978 331968 400046
rect 331648 399922 331718 399978
rect 331774 399922 331842 399978
rect 331898 399922 331968 399978
rect 331648 399888 331968 399922
rect 362368 400350 362688 400384
rect 362368 400294 362438 400350
rect 362494 400294 362562 400350
rect 362618 400294 362688 400350
rect 362368 400226 362688 400294
rect 362368 400170 362438 400226
rect 362494 400170 362562 400226
rect 362618 400170 362688 400226
rect 362368 400102 362688 400170
rect 362368 400046 362438 400102
rect 362494 400046 362562 400102
rect 362618 400046 362688 400102
rect 362368 399978 362688 400046
rect 362368 399922 362438 399978
rect 362494 399922 362562 399978
rect 362618 399922 362688 399978
rect 362368 399888 362688 399922
rect 393088 400350 393408 400384
rect 393088 400294 393158 400350
rect 393214 400294 393282 400350
rect 393338 400294 393408 400350
rect 393088 400226 393408 400294
rect 393088 400170 393158 400226
rect 393214 400170 393282 400226
rect 393338 400170 393408 400226
rect 393088 400102 393408 400170
rect 393088 400046 393158 400102
rect 393214 400046 393282 400102
rect 393338 400046 393408 400102
rect 393088 399978 393408 400046
rect 393088 399922 393158 399978
rect 393214 399922 393282 399978
rect 393338 399922 393408 399978
rect 393088 399888 393408 399922
rect 423808 400350 424128 400384
rect 423808 400294 423878 400350
rect 423934 400294 424002 400350
rect 424058 400294 424128 400350
rect 423808 400226 424128 400294
rect 423808 400170 423878 400226
rect 423934 400170 424002 400226
rect 424058 400170 424128 400226
rect 423808 400102 424128 400170
rect 423808 400046 423878 400102
rect 423934 400046 424002 400102
rect 424058 400046 424128 400102
rect 423808 399978 424128 400046
rect 423808 399922 423878 399978
rect 423934 399922 424002 399978
rect 424058 399922 424128 399978
rect 423808 399888 424128 399922
rect 454528 400350 454848 400384
rect 454528 400294 454598 400350
rect 454654 400294 454722 400350
rect 454778 400294 454848 400350
rect 454528 400226 454848 400294
rect 454528 400170 454598 400226
rect 454654 400170 454722 400226
rect 454778 400170 454848 400226
rect 454528 400102 454848 400170
rect 454528 400046 454598 400102
rect 454654 400046 454722 400102
rect 454778 400046 454848 400102
rect 454528 399978 454848 400046
rect 454528 399922 454598 399978
rect 454654 399922 454722 399978
rect 454778 399922 454848 399978
rect 454528 399888 454848 399922
rect 485248 400350 485568 400384
rect 485248 400294 485318 400350
rect 485374 400294 485442 400350
rect 485498 400294 485568 400350
rect 485248 400226 485568 400294
rect 485248 400170 485318 400226
rect 485374 400170 485442 400226
rect 485498 400170 485568 400226
rect 485248 400102 485568 400170
rect 485248 400046 485318 400102
rect 485374 400046 485442 400102
rect 485498 400046 485568 400102
rect 485248 399978 485568 400046
rect 485248 399922 485318 399978
rect 485374 399922 485442 399978
rect 485498 399922 485568 399978
rect 485248 399888 485568 399922
rect 515968 400350 516288 400384
rect 515968 400294 516038 400350
rect 516094 400294 516162 400350
rect 516218 400294 516288 400350
rect 515968 400226 516288 400294
rect 515968 400170 516038 400226
rect 516094 400170 516162 400226
rect 516218 400170 516288 400226
rect 515968 400102 516288 400170
rect 515968 400046 516038 400102
rect 516094 400046 516162 400102
rect 516218 400046 516288 400102
rect 515968 399978 516288 400046
rect 515968 399922 516038 399978
rect 516094 399922 516162 399978
rect 516218 399922 516288 399978
rect 515968 399888 516288 399922
rect 525154 400350 525774 417922
rect 525154 400294 525250 400350
rect 525306 400294 525374 400350
rect 525430 400294 525498 400350
rect 525554 400294 525622 400350
rect 525678 400294 525774 400350
rect 525154 400226 525774 400294
rect 525154 400170 525250 400226
rect 525306 400170 525374 400226
rect 525430 400170 525498 400226
rect 525554 400170 525622 400226
rect 525678 400170 525774 400226
rect 525154 400102 525774 400170
rect 525154 400046 525250 400102
rect 525306 400046 525374 400102
rect 525430 400046 525498 400102
rect 525554 400046 525622 400102
rect 525678 400046 525774 400102
rect 525154 399978 525774 400046
rect 525154 399922 525250 399978
rect 525306 399922 525374 399978
rect 525430 399922 525498 399978
rect 525554 399922 525622 399978
rect 525678 399922 525774 399978
rect 6874 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 7494 388350
rect 6874 388226 7494 388294
rect 6874 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 7494 388226
rect 6874 388102 7494 388170
rect 6874 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 7494 388102
rect 6874 387978 7494 388046
rect 6874 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 7494 387978
rect 6874 370350 7494 387922
rect 39808 388350 40128 388384
rect 39808 388294 39878 388350
rect 39934 388294 40002 388350
rect 40058 388294 40128 388350
rect 39808 388226 40128 388294
rect 39808 388170 39878 388226
rect 39934 388170 40002 388226
rect 40058 388170 40128 388226
rect 39808 388102 40128 388170
rect 39808 388046 39878 388102
rect 39934 388046 40002 388102
rect 40058 388046 40128 388102
rect 39808 387978 40128 388046
rect 39808 387922 39878 387978
rect 39934 387922 40002 387978
rect 40058 387922 40128 387978
rect 39808 387888 40128 387922
rect 70528 388350 70848 388384
rect 70528 388294 70598 388350
rect 70654 388294 70722 388350
rect 70778 388294 70848 388350
rect 70528 388226 70848 388294
rect 70528 388170 70598 388226
rect 70654 388170 70722 388226
rect 70778 388170 70848 388226
rect 70528 388102 70848 388170
rect 70528 388046 70598 388102
rect 70654 388046 70722 388102
rect 70778 388046 70848 388102
rect 70528 387978 70848 388046
rect 70528 387922 70598 387978
rect 70654 387922 70722 387978
rect 70778 387922 70848 387978
rect 70528 387888 70848 387922
rect 101248 388350 101568 388384
rect 101248 388294 101318 388350
rect 101374 388294 101442 388350
rect 101498 388294 101568 388350
rect 101248 388226 101568 388294
rect 101248 388170 101318 388226
rect 101374 388170 101442 388226
rect 101498 388170 101568 388226
rect 101248 388102 101568 388170
rect 101248 388046 101318 388102
rect 101374 388046 101442 388102
rect 101498 388046 101568 388102
rect 101248 387978 101568 388046
rect 101248 387922 101318 387978
rect 101374 387922 101442 387978
rect 101498 387922 101568 387978
rect 101248 387888 101568 387922
rect 131968 388350 132288 388384
rect 131968 388294 132038 388350
rect 132094 388294 132162 388350
rect 132218 388294 132288 388350
rect 131968 388226 132288 388294
rect 131968 388170 132038 388226
rect 132094 388170 132162 388226
rect 132218 388170 132288 388226
rect 131968 388102 132288 388170
rect 131968 388046 132038 388102
rect 132094 388046 132162 388102
rect 132218 388046 132288 388102
rect 131968 387978 132288 388046
rect 131968 387922 132038 387978
rect 132094 387922 132162 387978
rect 132218 387922 132288 387978
rect 131968 387888 132288 387922
rect 162688 388350 163008 388384
rect 162688 388294 162758 388350
rect 162814 388294 162882 388350
rect 162938 388294 163008 388350
rect 162688 388226 163008 388294
rect 162688 388170 162758 388226
rect 162814 388170 162882 388226
rect 162938 388170 163008 388226
rect 162688 388102 163008 388170
rect 162688 388046 162758 388102
rect 162814 388046 162882 388102
rect 162938 388046 163008 388102
rect 162688 387978 163008 388046
rect 162688 387922 162758 387978
rect 162814 387922 162882 387978
rect 162938 387922 163008 387978
rect 162688 387888 163008 387922
rect 193408 388350 193728 388384
rect 193408 388294 193478 388350
rect 193534 388294 193602 388350
rect 193658 388294 193728 388350
rect 193408 388226 193728 388294
rect 193408 388170 193478 388226
rect 193534 388170 193602 388226
rect 193658 388170 193728 388226
rect 193408 388102 193728 388170
rect 193408 388046 193478 388102
rect 193534 388046 193602 388102
rect 193658 388046 193728 388102
rect 193408 387978 193728 388046
rect 193408 387922 193478 387978
rect 193534 387922 193602 387978
rect 193658 387922 193728 387978
rect 193408 387888 193728 387922
rect 224128 388350 224448 388384
rect 224128 388294 224198 388350
rect 224254 388294 224322 388350
rect 224378 388294 224448 388350
rect 224128 388226 224448 388294
rect 224128 388170 224198 388226
rect 224254 388170 224322 388226
rect 224378 388170 224448 388226
rect 224128 388102 224448 388170
rect 224128 388046 224198 388102
rect 224254 388046 224322 388102
rect 224378 388046 224448 388102
rect 224128 387978 224448 388046
rect 224128 387922 224198 387978
rect 224254 387922 224322 387978
rect 224378 387922 224448 387978
rect 224128 387888 224448 387922
rect 254848 388350 255168 388384
rect 254848 388294 254918 388350
rect 254974 388294 255042 388350
rect 255098 388294 255168 388350
rect 254848 388226 255168 388294
rect 254848 388170 254918 388226
rect 254974 388170 255042 388226
rect 255098 388170 255168 388226
rect 254848 388102 255168 388170
rect 254848 388046 254918 388102
rect 254974 388046 255042 388102
rect 255098 388046 255168 388102
rect 254848 387978 255168 388046
rect 254848 387922 254918 387978
rect 254974 387922 255042 387978
rect 255098 387922 255168 387978
rect 254848 387888 255168 387922
rect 285568 388350 285888 388384
rect 285568 388294 285638 388350
rect 285694 388294 285762 388350
rect 285818 388294 285888 388350
rect 285568 388226 285888 388294
rect 285568 388170 285638 388226
rect 285694 388170 285762 388226
rect 285818 388170 285888 388226
rect 285568 388102 285888 388170
rect 285568 388046 285638 388102
rect 285694 388046 285762 388102
rect 285818 388046 285888 388102
rect 285568 387978 285888 388046
rect 285568 387922 285638 387978
rect 285694 387922 285762 387978
rect 285818 387922 285888 387978
rect 285568 387888 285888 387922
rect 316288 388350 316608 388384
rect 316288 388294 316358 388350
rect 316414 388294 316482 388350
rect 316538 388294 316608 388350
rect 316288 388226 316608 388294
rect 316288 388170 316358 388226
rect 316414 388170 316482 388226
rect 316538 388170 316608 388226
rect 316288 388102 316608 388170
rect 316288 388046 316358 388102
rect 316414 388046 316482 388102
rect 316538 388046 316608 388102
rect 316288 387978 316608 388046
rect 316288 387922 316358 387978
rect 316414 387922 316482 387978
rect 316538 387922 316608 387978
rect 316288 387888 316608 387922
rect 347008 388350 347328 388384
rect 347008 388294 347078 388350
rect 347134 388294 347202 388350
rect 347258 388294 347328 388350
rect 347008 388226 347328 388294
rect 347008 388170 347078 388226
rect 347134 388170 347202 388226
rect 347258 388170 347328 388226
rect 347008 388102 347328 388170
rect 347008 388046 347078 388102
rect 347134 388046 347202 388102
rect 347258 388046 347328 388102
rect 347008 387978 347328 388046
rect 347008 387922 347078 387978
rect 347134 387922 347202 387978
rect 347258 387922 347328 387978
rect 347008 387888 347328 387922
rect 377728 388350 378048 388384
rect 377728 388294 377798 388350
rect 377854 388294 377922 388350
rect 377978 388294 378048 388350
rect 377728 388226 378048 388294
rect 377728 388170 377798 388226
rect 377854 388170 377922 388226
rect 377978 388170 378048 388226
rect 377728 388102 378048 388170
rect 377728 388046 377798 388102
rect 377854 388046 377922 388102
rect 377978 388046 378048 388102
rect 377728 387978 378048 388046
rect 377728 387922 377798 387978
rect 377854 387922 377922 387978
rect 377978 387922 378048 387978
rect 377728 387888 378048 387922
rect 408448 388350 408768 388384
rect 408448 388294 408518 388350
rect 408574 388294 408642 388350
rect 408698 388294 408768 388350
rect 408448 388226 408768 388294
rect 408448 388170 408518 388226
rect 408574 388170 408642 388226
rect 408698 388170 408768 388226
rect 408448 388102 408768 388170
rect 408448 388046 408518 388102
rect 408574 388046 408642 388102
rect 408698 388046 408768 388102
rect 408448 387978 408768 388046
rect 408448 387922 408518 387978
rect 408574 387922 408642 387978
rect 408698 387922 408768 387978
rect 408448 387888 408768 387922
rect 439168 388350 439488 388384
rect 439168 388294 439238 388350
rect 439294 388294 439362 388350
rect 439418 388294 439488 388350
rect 439168 388226 439488 388294
rect 439168 388170 439238 388226
rect 439294 388170 439362 388226
rect 439418 388170 439488 388226
rect 439168 388102 439488 388170
rect 439168 388046 439238 388102
rect 439294 388046 439362 388102
rect 439418 388046 439488 388102
rect 439168 387978 439488 388046
rect 439168 387922 439238 387978
rect 439294 387922 439362 387978
rect 439418 387922 439488 387978
rect 439168 387888 439488 387922
rect 469888 388350 470208 388384
rect 469888 388294 469958 388350
rect 470014 388294 470082 388350
rect 470138 388294 470208 388350
rect 469888 388226 470208 388294
rect 469888 388170 469958 388226
rect 470014 388170 470082 388226
rect 470138 388170 470208 388226
rect 469888 388102 470208 388170
rect 469888 388046 469958 388102
rect 470014 388046 470082 388102
rect 470138 388046 470208 388102
rect 469888 387978 470208 388046
rect 469888 387922 469958 387978
rect 470014 387922 470082 387978
rect 470138 387922 470208 387978
rect 469888 387888 470208 387922
rect 500608 388350 500928 388384
rect 500608 388294 500678 388350
rect 500734 388294 500802 388350
rect 500858 388294 500928 388350
rect 500608 388226 500928 388294
rect 500608 388170 500678 388226
rect 500734 388170 500802 388226
rect 500858 388170 500928 388226
rect 500608 388102 500928 388170
rect 500608 388046 500678 388102
rect 500734 388046 500802 388102
rect 500858 388046 500928 388102
rect 500608 387978 500928 388046
rect 500608 387922 500678 387978
rect 500734 387922 500802 387978
rect 500858 387922 500928 387978
rect 500608 387888 500928 387922
rect 24448 382350 24768 382384
rect 24448 382294 24518 382350
rect 24574 382294 24642 382350
rect 24698 382294 24768 382350
rect 24448 382226 24768 382294
rect 24448 382170 24518 382226
rect 24574 382170 24642 382226
rect 24698 382170 24768 382226
rect 24448 382102 24768 382170
rect 24448 382046 24518 382102
rect 24574 382046 24642 382102
rect 24698 382046 24768 382102
rect 24448 381978 24768 382046
rect 24448 381922 24518 381978
rect 24574 381922 24642 381978
rect 24698 381922 24768 381978
rect 24448 381888 24768 381922
rect 55168 382350 55488 382384
rect 55168 382294 55238 382350
rect 55294 382294 55362 382350
rect 55418 382294 55488 382350
rect 55168 382226 55488 382294
rect 55168 382170 55238 382226
rect 55294 382170 55362 382226
rect 55418 382170 55488 382226
rect 55168 382102 55488 382170
rect 55168 382046 55238 382102
rect 55294 382046 55362 382102
rect 55418 382046 55488 382102
rect 55168 381978 55488 382046
rect 55168 381922 55238 381978
rect 55294 381922 55362 381978
rect 55418 381922 55488 381978
rect 55168 381888 55488 381922
rect 85888 382350 86208 382384
rect 85888 382294 85958 382350
rect 86014 382294 86082 382350
rect 86138 382294 86208 382350
rect 85888 382226 86208 382294
rect 85888 382170 85958 382226
rect 86014 382170 86082 382226
rect 86138 382170 86208 382226
rect 85888 382102 86208 382170
rect 85888 382046 85958 382102
rect 86014 382046 86082 382102
rect 86138 382046 86208 382102
rect 85888 381978 86208 382046
rect 85888 381922 85958 381978
rect 86014 381922 86082 381978
rect 86138 381922 86208 381978
rect 85888 381888 86208 381922
rect 116608 382350 116928 382384
rect 116608 382294 116678 382350
rect 116734 382294 116802 382350
rect 116858 382294 116928 382350
rect 116608 382226 116928 382294
rect 116608 382170 116678 382226
rect 116734 382170 116802 382226
rect 116858 382170 116928 382226
rect 116608 382102 116928 382170
rect 116608 382046 116678 382102
rect 116734 382046 116802 382102
rect 116858 382046 116928 382102
rect 116608 381978 116928 382046
rect 116608 381922 116678 381978
rect 116734 381922 116802 381978
rect 116858 381922 116928 381978
rect 116608 381888 116928 381922
rect 147328 382350 147648 382384
rect 147328 382294 147398 382350
rect 147454 382294 147522 382350
rect 147578 382294 147648 382350
rect 147328 382226 147648 382294
rect 147328 382170 147398 382226
rect 147454 382170 147522 382226
rect 147578 382170 147648 382226
rect 147328 382102 147648 382170
rect 147328 382046 147398 382102
rect 147454 382046 147522 382102
rect 147578 382046 147648 382102
rect 147328 381978 147648 382046
rect 147328 381922 147398 381978
rect 147454 381922 147522 381978
rect 147578 381922 147648 381978
rect 147328 381888 147648 381922
rect 178048 382350 178368 382384
rect 178048 382294 178118 382350
rect 178174 382294 178242 382350
rect 178298 382294 178368 382350
rect 178048 382226 178368 382294
rect 178048 382170 178118 382226
rect 178174 382170 178242 382226
rect 178298 382170 178368 382226
rect 178048 382102 178368 382170
rect 178048 382046 178118 382102
rect 178174 382046 178242 382102
rect 178298 382046 178368 382102
rect 178048 381978 178368 382046
rect 178048 381922 178118 381978
rect 178174 381922 178242 381978
rect 178298 381922 178368 381978
rect 178048 381888 178368 381922
rect 208768 382350 209088 382384
rect 208768 382294 208838 382350
rect 208894 382294 208962 382350
rect 209018 382294 209088 382350
rect 208768 382226 209088 382294
rect 208768 382170 208838 382226
rect 208894 382170 208962 382226
rect 209018 382170 209088 382226
rect 208768 382102 209088 382170
rect 208768 382046 208838 382102
rect 208894 382046 208962 382102
rect 209018 382046 209088 382102
rect 208768 381978 209088 382046
rect 208768 381922 208838 381978
rect 208894 381922 208962 381978
rect 209018 381922 209088 381978
rect 208768 381888 209088 381922
rect 239488 382350 239808 382384
rect 239488 382294 239558 382350
rect 239614 382294 239682 382350
rect 239738 382294 239808 382350
rect 239488 382226 239808 382294
rect 239488 382170 239558 382226
rect 239614 382170 239682 382226
rect 239738 382170 239808 382226
rect 239488 382102 239808 382170
rect 239488 382046 239558 382102
rect 239614 382046 239682 382102
rect 239738 382046 239808 382102
rect 239488 381978 239808 382046
rect 239488 381922 239558 381978
rect 239614 381922 239682 381978
rect 239738 381922 239808 381978
rect 239488 381888 239808 381922
rect 270208 382350 270528 382384
rect 270208 382294 270278 382350
rect 270334 382294 270402 382350
rect 270458 382294 270528 382350
rect 270208 382226 270528 382294
rect 270208 382170 270278 382226
rect 270334 382170 270402 382226
rect 270458 382170 270528 382226
rect 270208 382102 270528 382170
rect 270208 382046 270278 382102
rect 270334 382046 270402 382102
rect 270458 382046 270528 382102
rect 270208 381978 270528 382046
rect 270208 381922 270278 381978
rect 270334 381922 270402 381978
rect 270458 381922 270528 381978
rect 270208 381888 270528 381922
rect 300928 382350 301248 382384
rect 300928 382294 300998 382350
rect 301054 382294 301122 382350
rect 301178 382294 301248 382350
rect 300928 382226 301248 382294
rect 300928 382170 300998 382226
rect 301054 382170 301122 382226
rect 301178 382170 301248 382226
rect 300928 382102 301248 382170
rect 300928 382046 300998 382102
rect 301054 382046 301122 382102
rect 301178 382046 301248 382102
rect 300928 381978 301248 382046
rect 300928 381922 300998 381978
rect 301054 381922 301122 381978
rect 301178 381922 301248 381978
rect 300928 381888 301248 381922
rect 331648 382350 331968 382384
rect 331648 382294 331718 382350
rect 331774 382294 331842 382350
rect 331898 382294 331968 382350
rect 331648 382226 331968 382294
rect 331648 382170 331718 382226
rect 331774 382170 331842 382226
rect 331898 382170 331968 382226
rect 331648 382102 331968 382170
rect 331648 382046 331718 382102
rect 331774 382046 331842 382102
rect 331898 382046 331968 382102
rect 331648 381978 331968 382046
rect 331648 381922 331718 381978
rect 331774 381922 331842 381978
rect 331898 381922 331968 381978
rect 331648 381888 331968 381922
rect 362368 382350 362688 382384
rect 362368 382294 362438 382350
rect 362494 382294 362562 382350
rect 362618 382294 362688 382350
rect 362368 382226 362688 382294
rect 362368 382170 362438 382226
rect 362494 382170 362562 382226
rect 362618 382170 362688 382226
rect 362368 382102 362688 382170
rect 362368 382046 362438 382102
rect 362494 382046 362562 382102
rect 362618 382046 362688 382102
rect 362368 381978 362688 382046
rect 362368 381922 362438 381978
rect 362494 381922 362562 381978
rect 362618 381922 362688 381978
rect 362368 381888 362688 381922
rect 393088 382350 393408 382384
rect 393088 382294 393158 382350
rect 393214 382294 393282 382350
rect 393338 382294 393408 382350
rect 393088 382226 393408 382294
rect 393088 382170 393158 382226
rect 393214 382170 393282 382226
rect 393338 382170 393408 382226
rect 393088 382102 393408 382170
rect 393088 382046 393158 382102
rect 393214 382046 393282 382102
rect 393338 382046 393408 382102
rect 393088 381978 393408 382046
rect 393088 381922 393158 381978
rect 393214 381922 393282 381978
rect 393338 381922 393408 381978
rect 393088 381888 393408 381922
rect 423808 382350 424128 382384
rect 423808 382294 423878 382350
rect 423934 382294 424002 382350
rect 424058 382294 424128 382350
rect 423808 382226 424128 382294
rect 423808 382170 423878 382226
rect 423934 382170 424002 382226
rect 424058 382170 424128 382226
rect 423808 382102 424128 382170
rect 423808 382046 423878 382102
rect 423934 382046 424002 382102
rect 424058 382046 424128 382102
rect 423808 381978 424128 382046
rect 423808 381922 423878 381978
rect 423934 381922 424002 381978
rect 424058 381922 424128 381978
rect 423808 381888 424128 381922
rect 454528 382350 454848 382384
rect 454528 382294 454598 382350
rect 454654 382294 454722 382350
rect 454778 382294 454848 382350
rect 454528 382226 454848 382294
rect 454528 382170 454598 382226
rect 454654 382170 454722 382226
rect 454778 382170 454848 382226
rect 454528 382102 454848 382170
rect 454528 382046 454598 382102
rect 454654 382046 454722 382102
rect 454778 382046 454848 382102
rect 454528 381978 454848 382046
rect 454528 381922 454598 381978
rect 454654 381922 454722 381978
rect 454778 381922 454848 381978
rect 454528 381888 454848 381922
rect 485248 382350 485568 382384
rect 485248 382294 485318 382350
rect 485374 382294 485442 382350
rect 485498 382294 485568 382350
rect 485248 382226 485568 382294
rect 485248 382170 485318 382226
rect 485374 382170 485442 382226
rect 485498 382170 485568 382226
rect 485248 382102 485568 382170
rect 485248 382046 485318 382102
rect 485374 382046 485442 382102
rect 485498 382046 485568 382102
rect 485248 381978 485568 382046
rect 485248 381922 485318 381978
rect 485374 381922 485442 381978
rect 485498 381922 485568 381978
rect 485248 381888 485568 381922
rect 515968 382350 516288 382384
rect 515968 382294 516038 382350
rect 516094 382294 516162 382350
rect 516218 382294 516288 382350
rect 515968 382226 516288 382294
rect 515968 382170 516038 382226
rect 516094 382170 516162 382226
rect 516218 382170 516288 382226
rect 515968 382102 516288 382170
rect 515968 382046 516038 382102
rect 516094 382046 516162 382102
rect 516218 382046 516288 382102
rect 515968 381978 516288 382046
rect 515968 381922 516038 381978
rect 516094 381922 516162 381978
rect 516218 381922 516288 381978
rect 515968 381888 516288 381922
rect 525154 382350 525774 399922
rect 525154 382294 525250 382350
rect 525306 382294 525374 382350
rect 525430 382294 525498 382350
rect 525554 382294 525622 382350
rect 525678 382294 525774 382350
rect 525154 382226 525774 382294
rect 525154 382170 525250 382226
rect 525306 382170 525374 382226
rect 525430 382170 525498 382226
rect 525554 382170 525622 382226
rect 525678 382170 525774 382226
rect 525154 382102 525774 382170
rect 525154 382046 525250 382102
rect 525306 382046 525374 382102
rect 525430 382046 525498 382102
rect 525554 382046 525622 382102
rect 525678 382046 525774 382102
rect 525154 381978 525774 382046
rect 525154 381922 525250 381978
rect 525306 381922 525374 381978
rect 525430 381922 525498 381978
rect 525554 381922 525622 381978
rect 525678 381922 525774 381978
rect 6874 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 7494 370350
rect 6874 370226 7494 370294
rect 6874 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 7494 370226
rect 6874 370102 7494 370170
rect 6874 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 7494 370102
rect 6874 369978 7494 370046
rect 6874 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 7494 369978
rect 6874 352350 7494 369922
rect 39808 370350 40128 370384
rect 39808 370294 39878 370350
rect 39934 370294 40002 370350
rect 40058 370294 40128 370350
rect 39808 370226 40128 370294
rect 39808 370170 39878 370226
rect 39934 370170 40002 370226
rect 40058 370170 40128 370226
rect 39808 370102 40128 370170
rect 39808 370046 39878 370102
rect 39934 370046 40002 370102
rect 40058 370046 40128 370102
rect 39808 369978 40128 370046
rect 39808 369922 39878 369978
rect 39934 369922 40002 369978
rect 40058 369922 40128 369978
rect 39808 369888 40128 369922
rect 70528 370350 70848 370384
rect 70528 370294 70598 370350
rect 70654 370294 70722 370350
rect 70778 370294 70848 370350
rect 70528 370226 70848 370294
rect 70528 370170 70598 370226
rect 70654 370170 70722 370226
rect 70778 370170 70848 370226
rect 70528 370102 70848 370170
rect 70528 370046 70598 370102
rect 70654 370046 70722 370102
rect 70778 370046 70848 370102
rect 70528 369978 70848 370046
rect 70528 369922 70598 369978
rect 70654 369922 70722 369978
rect 70778 369922 70848 369978
rect 70528 369888 70848 369922
rect 101248 370350 101568 370384
rect 101248 370294 101318 370350
rect 101374 370294 101442 370350
rect 101498 370294 101568 370350
rect 101248 370226 101568 370294
rect 101248 370170 101318 370226
rect 101374 370170 101442 370226
rect 101498 370170 101568 370226
rect 101248 370102 101568 370170
rect 101248 370046 101318 370102
rect 101374 370046 101442 370102
rect 101498 370046 101568 370102
rect 101248 369978 101568 370046
rect 101248 369922 101318 369978
rect 101374 369922 101442 369978
rect 101498 369922 101568 369978
rect 101248 369888 101568 369922
rect 131968 370350 132288 370384
rect 131968 370294 132038 370350
rect 132094 370294 132162 370350
rect 132218 370294 132288 370350
rect 131968 370226 132288 370294
rect 131968 370170 132038 370226
rect 132094 370170 132162 370226
rect 132218 370170 132288 370226
rect 131968 370102 132288 370170
rect 131968 370046 132038 370102
rect 132094 370046 132162 370102
rect 132218 370046 132288 370102
rect 131968 369978 132288 370046
rect 131968 369922 132038 369978
rect 132094 369922 132162 369978
rect 132218 369922 132288 369978
rect 131968 369888 132288 369922
rect 162688 370350 163008 370384
rect 162688 370294 162758 370350
rect 162814 370294 162882 370350
rect 162938 370294 163008 370350
rect 162688 370226 163008 370294
rect 162688 370170 162758 370226
rect 162814 370170 162882 370226
rect 162938 370170 163008 370226
rect 162688 370102 163008 370170
rect 162688 370046 162758 370102
rect 162814 370046 162882 370102
rect 162938 370046 163008 370102
rect 162688 369978 163008 370046
rect 162688 369922 162758 369978
rect 162814 369922 162882 369978
rect 162938 369922 163008 369978
rect 162688 369888 163008 369922
rect 193408 370350 193728 370384
rect 193408 370294 193478 370350
rect 193534 370294 193602 370350
rect 193658 370294 193728 370350
rect 193408 370226 193728 370294
rect 193408 370170 193478 370226
rect 193534 370170 193602 370226
rect 193658 370170 193728 370226
rect 193408 370102 193728 370170
rect 193408 370046 193478 370102
rect 193534 370046 193602 370102
rect 193658 370046 193728 370102
rect 193408 369978 193728 370046
rect 193408 369922 193478 369978
rect 193534 369922 193602 369978
rect 193658 369922 193728 369978
rect 193408 369888 193728 369922
rect 224128 370350 224448 370384
rect 224128 370294 224198 370350
rect 224254 370294 224322 370350
rect 224378 370294 224448 370350
rect 224128 370226 224448 370294
rect 224128 370170 224198 370226
rect 224254 370170 224322 370226
rect 224378 370170 224448 370226
rect 224128 370102 224448 370170
rect 224128 370046 224198 370102
rect 224254 370046 224322 370102
rect 224378 370046 224448 370102
rect 224128 369978 224448 370046
rect 224128 369922 224198 369978
rect 224254 369922 224322 369978
rect 224378 369922 224448 369978
rect 224128 369888 224448 369922
rect 254848 370350 255168 370384
rect 254848 370294 254918 370350
rect 254974 370294 255042 370350
rect 255098 370294 255168 370350
rect 254848 370226 255168 370294
rect 254848 370170 254918 370226
rect 254974 370170 255042 370226
rect 255098 370170 255168 370226
rect 254848 370102 255168 370170
rect 254848 370046 254918 370102
rect 254974 370046 255042 370102
rect 255098 370046 255168 370102
rect 254848 369978 255168 370046
rect 254848 369922 254918 369978
rect 254974 369922 255042 369978
rect 255098 369922 255168 369978
rect 254848 369888 255168 369922
rect 285568 370350 285888 370384
rect 285568 370294 285638 370350
rect 285694 370294 285762 370350
rect 285818 370294 285888 370350
rect 285568 370226 285888 370294
rect 285568 370170 285638 370226
rect 285694 370170 285762 370226
rect 285818 370170 285888 370226
rect 285568 370102 285888 370170
rect 285568 370046 285638 370102
rect 285694 370046 285762 370102
rect 285818 370046 285888 370102
rect 285568 369978 285888 370046
rect 285568 369922 285638 369978
rect 285694 369922 285762 369978
rect 285818 369922 285888 369978
rect 285568 369888 285888 369922
rect 316288 370350 316608 370384
rect 316288 370294 316358 370350
rect 316414 370294 316482 370350
rect 316538 370294 316608 370350
rect 316288 370226 316608 370294
rect 316288 370170 316358 370226
rect 316414 370170 316482 370226
rect 316538 370170 316608 370226
rect 316288 370102 316608 370170
rect 316288 370046 316358 370102
rect 316414 370046 316482 370102
rect 316538 370046 316608 370102
rect 316288 369978 316608 370046
rect 316288 369922 316358 369978
rect 316414 369922 316482 369978
rect 316538 369922 316608 369978
rect 316288 369888 316608 369922
rect 347008 370350 347328 370384
rect 347008 370294 347078 370350
rect 347134 370294 347202 370350
rect 347258 370294 347328 370350
rect 347008 370226 347328 370294
rect 347008 370170 347078 370226
rect 347134 370170 347202 370226
rect 347258 370170 347328 370226
rect 347008 370102 347328 370170
rect 347008 370046 347078 370102
rect 347134 370046 347202 370102
rect 347258 370046 347328 370102
rect 347008 369978 347328 370046
rect 347008 369922 347078 369978
rect 347134 369922 347202 369978
rect 347258 369922 347328 369978
rect 347008 369888 347328 369922
rect 377728 370350 378048 370384
rect 377728 370294 377798 370350
rect 377854 370294 377922 370350
rect 377978 370294 378048 370350
rect 377728 370226 378048 370294
rect 377728 370170 377798 370226
rect 377854 370170 377922 370226
rect 377978 370170 378048 370226
rect 377728 370102 378048 370170
rect 377728 370046 377798 370102
rect 377854 370046 377922 370102
rect 377978 370046 378048 370102
rect 377728 369978 378048 370046
rect 377728 369922 377798 369978
rect 377854 369922 377922 369978
rect 377978 369922 378048 369978
rect 377728 369888 378048 369922
rect 408448 370350 408768 370384
rect 408448 370294 408518 370350
rect 408574 370294 408642 370350
rect 408698 370294 408768 370350
rect 408448 370226 408768 370294
rect 408448 370170 408518 370226
rect 408574 370170 408642 370226
rect 408698 370170 408768 370226
rect 408448 370102 408768 370170
rect 408448 370046 408518 370102
rect 408574 370046 408642 370102
rect 408698 370046 408768 370102
rect 408448 369978 408768 370046
rect 408448 369922 408518 369978
rect 408574 369922 408642 369978
rect 408698 369922 408768 369978
rect 408448 369888 408768 369922
rect 439168 370350 439488 370384
rect 439168 370294 439238 370350
rect 439294 370294 439362 370350
rect 439418 370294 439488 370350
rect 439168 370226 439488 370294
rect 439168 370170 439238 370226
rect 439294 370170 439362 370226
rect 439418 370170 439488 370226
rect 439168 370102 439488 370170
rect 439168 370046 439238 370102
rect 439294 370046 439362 370102
rect 439418 370046 439488 370102
rect 439168 369978 439488 370046
rect 439168 369922 439238 369978
rect 439294 369922 439362 369978
rect 439418 369922 439488 369978
rect 439168 369888 439488 369922
rect 469888 370350 470208 370384
rect 469888 370294 469958 370350
rect 470014 370294 470082 370350
rect 470138 370294 470208 370350
rect 469888 370226 470208 370294
rect 469888 370170 469958 370226
rect 470014 370170 470082 370226
rect 470138 370170 470208 370226
rect 469888 370102 470208 370170
rect 469888 370046 469958 370102
rect 470014 370046 470082 370102
rect 470138 370046 470208 370102
rect 469888 369978 470208 370046
rect 469888 369922 469958 369978
rect 470014 369922 470082 369978
rect 470138 369922 470208 369978
rect 469888 369888 470208 369922
rect 500608 370350 500928 370384
rect 500608 370294 500678 370350
rect 500734 370294 500802 370350
rect 500858 370294 500928 370350
rect 500608 370226 500928 370294
rect 500608 370170 500678 370226
rect 500734 370170 500802 370226
rect 500858 370170 500928 370226
rect 500608 370102 500928 370170
rect 500608 370046 500678 370102
rect 500734 370046 500802 370102
rect 500858 370046 500928 370102
rect 500608 369978 500928 370046
rect 500608 369922 500678 369978
rect 500734 369922 500802 369978
rect 500858 369922 500928 369978
rect 500608 369888 500928 369922
rect 24448 364350 24768 364384
rect 24448 364294 24518 364350
rect 24574 364294 24642 364350
rect 24698 364294 24768 364350
rect 24448 364226 24768 364294
rect 24448 364170 24518 364226
rect 24574 364170 24642 364226
rect 24698 364170 24768 364226
rect 24448 364102 24768 364170
rect 24448 364046 24518 364102
rect 24574 364046 24642 364102
rect 24698 364046 24768 364102
rect 24448 363978 24768 364046
rect 24448 363922 24518 363978
rect 24574 363922 24642 363978
rect 24698 363922 24768 363978
rect 24448 363888 24768 363922
rect 55168 364350 55488 364384
rect 55168 364294 55238 364350
rect 55294 364294 55362 364350
rect 55418 364294 55488 364350
rect 55168 364226 55488 364294
rect 55168 364170 55238 364226
rect 55294 364170 55362 364226
rect 55418 364170 55488 364226
rect 55168 364102 55488 364170
rect 55168 364046 55238 364102
rect 55294 364046 55362 364102
rect 55418 364046 55488 364102
rect 55168 363978 55488 364046
rect 55168 363922 55238 363978
rect 55294 363922 55362 363978
rect 55418 363922 55488 363978
rect 55168 363888 55488 363922
rect 85888 364350 86208 364384
rect 85888 364294 85958 364350
rect 86014 364294 86082 364350
rect 86138 364294 86208 364350
rect 85888 364226 86208 364294
rect 85888 364170 85958 364226
rect 86014 364170 86082 364226
rect 86138 364170 86208 364226
rect 85888 364102 86208 364170
rect 85888 364046 85958 364102
rect 86014 364046 86082 364102
rect 86138 364046 86208 364102
rect 85888 363978 86208 364046
rect 85888 363922 85958 363978
rect 86014 363922 86082 363978
rect 86138 363922 86208 363978
rect 85888 363888 86208 363922
rect 116608 364350 116928 364384
rect 116608 364294 116678 364350
rect 116734 364294 116802 364350
rect 116858 364294 116928 364350
rect 116608 364226 116928 364294
rect 116608 364170 116678 364226
rect 116734 364170 116802 364226
rect 116858 364170 116928 364226
rect 116608 364102 116928 364170
rect 116608 364046 116678 364102
rect 116734 364046 116802 364102
rect 116858 364046 116928 364102
rect 116608 363978 116928 364046
rect 116608 363922 116678 363978
rect 116734 363922 116802 363978
rect 116858 363922 116928 363978
rect 116608 363888 116928 363922
rect 147328 364350 147648 364384
rect 147328 364294 147398 364350
rect 147454 364294 147522 364350
rect 147578 364294 147648 364350
rect 147328 364226 147648 364294
rect 147328 364170 147398 364226
rect 147454 364170 147522 364226
rect 147578 364170 147648 364226
rect 147328 364102 147648 364170
rect 147328 364046 147398 364102
rect 147454 364046 147522 364102
rect 147578 364046 147648 364102
rect 147328 363978 147648 364046
rect 147328 363922 147398 363978
rect 147454 363922 147522 363978
rect 147578 363922 147648 363978
rect 147328 363888 147648 363922
rect 178048 364350 178368 364384
rect 178048 364294 178118 364350
rect 178174 364294 178242 364350
rect 178298 364294 178368 364350
rect 178048 364226 178368 364294
rect 178048 364170 178118 364226
rect 178174 364170 178242 364226
rect 178298 364170 178368 364226
rect 178048 364102 178368 364170
rect 178048 364046 178118 364102
rect 178174 364046 178242 364102
rect 178298 364046 178368 364102
rect 178048 363978 178368 364046
rect 178048 363922 178118 363978
rect 178174 363922 178242 363978
rect 178298 363922 178368 363978
rect 178048 363888 178368 363922
rect 208768 364350 209088 364384
rect 208768 364294 208838 364350
rect 208894 364294 208962 364350
rect 209018 364294 209088 364350
rect 208768 364226 209088 364294
rect 208768 364170 208838 364226
rect 208894 364170 208962 364226
rect 209018 364170 209088 364226
rect 208768 364102 209088 364170
rect 208768 364046 208838 364102
rect 208894 364046 208962 364102
rect 209018 364046 209088 364102
rect 208768 363978 209088 364046
rect 208768 363922 208838 363978
rect 208894 363922 208962 363978
rect 209018 363922 209088 363978
rect 208768 363888 209088 363922
rect 239488 364350 239808 364384
rect 239488 364294 239558 364350
rect 239614 364294 239682 364350
rect 239738 364294 239808 364350
rect 239488 364226 239808 364294
rect 239488 364170 239558 364226
rect 239614 364170 239682 364226
rect 239738 364170 239808 364226
rect 239488 364102 239808 364170
rect 239488 364046 239558 364102
rect 239614 364046 239682 364102
rect 239738 364046 239808 364102
rect 239488 363978 239808 364046
rect 239488 363922 239558 363978
rect 239614 363922 239682 363978
rect 239738 363922 239808 363978
rect 239488 363888 239808 363922
rect 270208 364350 270528 364384
rect 270208 364294 270278 364350
rect 270334 364294 270402 364350
rect 270458 364294 270528 364350
rect 270208 364226 270528 364294
rect 270208 364170 270278 364226
rect 270334 364170 270402 364226
rect 270458 364170 270528 364226
rect 270208 364102 270528 364170
rect 270208 364046 270278 364102
rect 270334 364046 270402 364102
rect 270458 364046 270528 364102
rect 270208 363978 270528 364046
rect 270208 363922 270278 363978
rect 270334 363922 270402 363978
rect 270458 363922 270528 363978
rect 270208 363888 270528 363922
rect 300928 364350 301248 364384
rect 300928 364294 300998 364350
rect 301054 364294 301122 364350
rect 301178 364294 301248 364350
rect 300928 364226 301248 364294
rect 300928 364170 300998 364226
rect 301054 364170 301122 364226
rect 301178 364170 301248 364226
rect 300928 364102 301248 364170
rect 300928 364046 300998 364102
rect 301054 364046 301122 364102
rect 301178 364046 301248 364102
rect 300928 363978 301248 364046
rect 300928 363922 300998 363978
rect 301054 363922 301122 363978
rect 301178 363922 301248 363978
rect 300928 363888 301248 363922
rect 331648 364350 331968 364384
rect 331648 364294 331718 364350
rect 331774 364294 331842 364350
rect 331898 364294 331968 364350
rect 331648 364226 331968 364294
rect 331648 364170 331718 364226
rect 331774 364170 331842 364226
rect 331898 364170 331968 364226
rect 331648 364102 331968 364170
rect 331648 364046 331718 364102
rect 331774 364046 331842 364102
rect 331898 364046 331968 364102
rect 331648 363978 331968 364046
rect 331648 363922 331718 363978
rect 331774 363922 331842 363978
rect 331898 363922 331968 363978
rect 331648 363888 331968 363922
rect 362368 364350 362688 364384
rect 362368 364294 362438 364350
rect 362494 364294 362562 364350
rect 362618 364294 362688 364350
rect 362368 364226 362688 364294
rect 362368 364170 362438 364226
rect 362494 364170 362562 364226
rect 362618 364170 362688 364226
rect 362368 364102 362688 364170
rect 362368 364046 362438 364102
rect 362494 364046 362562 364102
rect 362618 364046 362688 364102
rect 362368 363978 362688 364046
rect 362368 363922 362438 363978
rect 362494 363922 362562 363978
rect 362618 363922 362688 363978
rect 362368 363888 362688 363922
rect 393088 364350 393408 364384
rect 393088 364294 393158 364350
rect 393214 364294 393282 364350
rect 393338 364294 393408 364350
rect 393088 364226 393408 364294
rect 393088 364170 393158 364226
rect 393214 364170 393282 364226
rect 393338 364170 393408 364226
rect 393088 364102 393408 364170
rect 393088 364046 393158 364102
rect 393214 364046 393282 364102
rect 393338 364046 393408 364102
rect 393088 363978 393408 364046
rect 393088 363922 393158 363978
rect 393214 363922 393282 363978
rect 393338 363922 393408 363978
rect 393088 363888 393408 363922
rect 423808 364350 424128 364384
rect 423808 364294 423878 364350
rect 423934 364294 424002 364350
rect 424058 364294 424128 364350
rect 423808 364226 424128 364294
rect 423808 364170 423878 364226
rect 423934 364170 424002 364226
rect 424058 364170 424128 364226
rect 423808 364102 424128 364170
rect 423808 364046 423878 364102
rect 423934 364046 424002 364102
rect 424058 364046 424128 364102
rect 423808 363978 424128 364046
rect 423808 363922 423878 363978
rect 423934 363922 424002 363978
rect 424058 363922 424128 363978
rect 423808 363888 424128 363922
rect 454528 364350 454848 364384
rect 454528 364294 454598 364350
rect 454654 364294 454722 364350
rect 454778 364294 454848 364350
rect 454528 364226 454848 364294
rect 454528 364170 454598 364226
rect 454654 364170 454722 364226
rect 454778 364170 454848 364226
rect 454528 364102 454848 364170
rect 454528 364046 454598 364102
rect 454654 364046 454722 364102
rect 454778 364046 454848 364102
rect 454528 363978 454848 364046
rect 454528 363922 454598 363978
rect 454654 363922 454722 363978
rect 454778 363922 454848 363978
rect 454528 363888 454848 363922
rect 485248 364350 485568 364384
rect 485248 364294 485318 364350
rect 485374 364294 485442 364350
rect 485498 364294 485568 364350
rect 485248 364226 485568 364294
rect 485248 364170 485318 364226
rect 485374 364170 485442 364226
rect 485498 364170 485568 364226
rect 485248 364102 485568 364170
rect 485248 364046 485318 364102
rect 485374 364046 485442 364102
rect 485498 364046 485568 364102
rect 485248 363978 485568 364046
rect 485248 363922 485318 363978
rect 485374 363922 485442 363978
rect 485498 363922 485568 363978
rect 485248 363888 485568 363922
rect 515968 364350 516288 364384
rect 515968 364294 516038 364350
rect 516094 364294 516162 364350
rect 516218 364294 516288 364350
rect 515968 364226 516288 364294
rect 515968 364170 516038 364226
rect 516094 364170 516162 364226
rect 516218 364170 516288 364226
rect 515968 364102 516288 364170
rect 515968 364046 516038 364102
rect 516094 364046 516162 364102
rect 516218 364046 516288 364102
rect 515968 363978 516288 364046
rect 515968 363922 516038 363978
rect 516094 363922 516162 363978
rect 516218 363922 516288 363978
rect 515968 363888 516288 363922
rect 525154 364350 525774 381922
rect 525154 364294 525250 364350
rect 525306 364294 525374 364350
rect 525430 364294 525498 364350
rect 525554 364294 525622 364350
rect 525678 364294 525774 364350
rect 525154 364226 525774 364294
rect 525154 364170 525250 364226
rect 525306 364170 525374 364226
rect 525430 364170 525498 364226
rect 525554 364170 525622 364226
rect 525678 364170 525774 364226
rect 525154 364102 525774 364170
rect 525154 364046 525250 364102
rect 525306 364046 525374 364102
rect 525430 364046 525498 364102
rect 525554 364046 525622 364102
rect 525678 364046 525774 364102
rect 525154 363978 525774 364046
rect 525154 363922 525250 363978
rect 525306 363922 525374 363978
rect 525430 363922 525498 363978
rect 525554 363922 525622 363978
rect 525678 363922 525774 363978
rect 6874 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 7494 352350
rect 6874 352226 7494 352294
rect 6874 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 7494 352226
rect 6874 352102 7494 352170
rect 6874 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 7494 352102
rect 6874 351978 7494 352046
rect 6874 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 7494 351978
rect 6874 334350 7494 351922
rect 39808 352350 40128 352384
rect 39808 352294 39878 352350
rect 39934 352294 40002 352350
rect 40058 352294 40128 352350
rect 39808 352226 40128 352294
rect 39808 352170 39878 352226
rect 39934 352170 40002 352226
rect 40058 352170 40128 352226
rect 39808 352102 40128 352170
rect 39808 352046 39878 352102
rect 39934 352046 40002 352102
rect 40058 352046 40128 352102
rect 39808 351978 40128 352046
rect 39808 351922 39878 351978
rect 39934 351922 40002 351978
rect 40058 351922 40128 351978
rect 39808 351888 40128 351922
rect 70528 352350 70848 352384
rect 70528 352294 70598 352350
rect 70654 352294 70722 352350
rect 70778 352294 70848 352350
rect 70528 352226 70848 352294
rect 70528 352170 70598 352226
rect 70654 352170 70722 352226
rect 70778 352170 70848 352226
rect 70528 352102 70848 352170
rect 70528 352046 70598 352102
rect 70654 352046 70722 352102
rect 70778 352046 70848 352102
rect 70528 351978 70848 352046
rect 70528 351922 70598 351978
rect 70654 351922 70722 351978
rect 70778 351922 70848 351978
rect 70528 351888 70848 351922
rect 101248 352350 101568 352384
rect 101248 352294 101318 352350
rect 101374 352294 101442 352350
rect 101498 352294 101568 352350
rect 101248 352226 101568 352294
rect 101248 352170 101318 352226
rect 101374 352170 101442 352226
rect 101498 352170 101568 352226
rect 101248 352102 101568 352170
rect 101248 352046 101318 352102
rect 101374 352046 101442 352102
rect 101498 352046 101568 352102
rect 101248 351978 101568 352046
rect 101248 351922 101318 351978
rect 101374 351922 101442 351978
rect 101498 351922 101568 351978
rect 101248 351888 101568 351922
rect 131968 352350 132288 352384
rect 131968 352294 132038 352350
rect 132094 352294 132162 352350
rect 132218 352294 132288 352350
rect 131968 352226 132288 352294
rect 131968 352170 132038 352226
rect 132094 352170 132162 352226
rect 132218 352170 132288 352226
rect 131968 352102 132288 352170
rect 131968 352046 132038 352102
rect 132094 352046 132162 352102
rect 132218 352046 132288 352102
rect 131968 351978 132288 352046
rect 131968 351922 132038 351978
rect 132094 351922 132162 351978
rect 132218 351922 132288 351978
rect 131968 351888 132288 351922
rect 162688 352350 163008 352384
rect 162688 352294 162758 352350
rect 162814 352294 162882 352350
rect 162938 352294 163008 352350
rect 162688 352226 163008 352294
rect 162688 352170 162758 352226
rect 162814 352170 162882 352226
rect 162938 352170 163008 352226
rect 162688 352102 163008 352170
rect 162688 352046 162758 352102
rect 162814 352046 162882 352102
rect 162938 352046 163008 352102
rect 162688 351978 163008 352046
rect 162688 351922 162758 351978
rect 162814 351922 162882 351978
rect 162938 351922 163008 351978
rect 162688 351888 163008 351922
rect 193408 352350 193728 352384
rect 193408 352294 193478 352350
rect 193534 352294 193602 352350
rect 193658 352294 193728 352350
rect 193408 352226 193728 352294
rect 193408 352170 193478 352226
rect 193534 352170 193602 352226
rect 193658 352170 193728 352226
rect 193408 352102 193728 352170
rect 193408 352046 193478 352102
rect 193534 352046 193602 352102
rect 193658 352046 193728 352102
rect 193408 351978 193728 352046
rect 193408 351922 193478 351978
rect 193534 351922 193602 351978
rect 193658 351922 193728 351978
rect 193408 351888 193728 351922
rect 224128 352350 224448 352384
rect 224128 352294 224198 352350
rect 224254 352294 224322 352350
rect 224378 352294 224448 352350
rect 224128 352226 224448 352294
rect 224128 352170 224198 352226
rect 224254 352170 224322 352226
rect 224378 352170 224448 352226
rect 224128 352102 224448 352170
rect 224128 352046 224198 352102
rect 224254 352046 224322 352102
rect 224378 352046 224448 352102
rect 224128 351978 224448 352046
rect 224128 351922 224198 351978
rect 224254 351922 224322 351978
rect 224378 351922 224448 351978
rect 224128 351888 224448 351922
rect 254848 352350 255168 352384
rect 254848 352294 254918 352350
rect 254974 352294 255042 352350
rect 255098 352294 255168 352350
rect 254848 352226 255168 352294
rect 254848 352170 254918 352226
rect 254974 352170 255042 352226
rect 255098 352170 255168 352226
rect 254848 352102 255168 352170
rect 254848 352046 254918 352102
rect 254974 352046 255042 352102
rect 255098 352046 255168 352102
rect 254848 351978 255168 352046
rect 254848 351922 254918 351978
rect 254974 351922 255042 351978
rect 255098 351922 255168 351978
rect 254848 351888 255168 351922
rect 285568 352350 285888 352384
rect 285568 352294 285638 352350
rect 285694 352294 285762 352350
rect 285818 352294 285888 352350
rect 285568 352226 285888 352294
rect 285568 352170 285638 352226
rect 285694 352170 285762 352226
rect 285818 352170 285888 352226
rect 285568 352102 285888 352170
rect 285568 352046 285638 352102
rect 285694 352046 285762 352102
rect 285818 352046 285888 352102
rect 285568 351978 285888 352046
rect 285568 351922 285638 351978
rect 285694 351922 285762 351978
rect 285818 351922 285888 351978
rect 285568 351888 285888 351922
rect 316288 352350 316608 352384
rect 316288 352294 316358 352350
rect 316414 352294 316482 352350
rect 316538 352294 316608 352350
rect 316288 352226 316608 352294
rect 316288 352170 316358 352226
rect 316414 352170 316482 352226
rect 316538 352170 316608 352226
rect 316288 352102 316608 352170
rect 316288 352046 316358 352102
rect 316414 352046 316482 352102
rect 316538 352046 316608 352102
rect 316288 351978 316608 352046
rect 316288 351922 316358 351978
rect 316414 351922 316482 351978
rect 316538 351922 316608 351978
rect 316288 351888 316608 351922
rect 347008 352350 347328 352384
rect 347008 352294 347078 352350
rect 347134 352294 347202 352350
rect 347258 352294 347328 352350
rect 347008 352226 347328 352294
rect 347008 352170 347078 352226
rect 347134 352170 347202 352226
rect 347258 352170 347328 352226
rect 347008 352102 347328 352170
rect 347008 352046 347078 352102
rect 347134 352046 347202 352102
rect 347258 352046 347328 352102
rect 347008 351978 347328 352046
rect 347008 351922 347078 351978
rect 347134 351922 347202 351978
rect 347258 351922 347328 351978
rect 347008 351888 347328 351922
rect 377728 352350 378048 352384
rect 377728 352294 377798 352350
rect 377854 352294 377922 352350
rect 377978 352294 378048 352350
rect 377728 352226 378048 352294
rect 377728 352170 377798 352226
rect 377854 352170 377922 352226
rect 377978 352170 378048 352226
rect 377728 352102 378048 352170
rect 377728 352046 377798 352102
rect 377854 352046 377922 352102
rect 377978 352046 378048 352102
rect 377728 351978 378048 352046
rect 377728 351922 377798 351978
rect 377854 351922 377922 351978
rect 377978 351922 378048 351978
rect 377728 351888 378048 351922
rect 408448 352350 408768 352384
rect 408448 352294 408518 352350
rect 408574 352294 408642 352350
rect 408698 352294 408768 352350
rect 408448 352226 408768 352294
rect 408448 352170 408518 352226
rect 408574 352170 408642 352226
rect 408698 352170 408768 352226
rect 408448 352102 408768 352170
rect 408448 352046 408518 352102
rect 408574 352046 408642 352102
rect 408698 352046 408768 352102
rect 408448 351978 408768 352046
rect 408448 351922 408518 351978
rect 408574 351922 408642 351978
rect 408698 351922 408768 351978
rect 408448 351888 408768 351922
rect 439168 352350 439488 352384
rect 439168 352294 439238 352350
rect 439294 352294 439362 352350
rect 439418 352294 439488 352350
rect 439168 352226 439488 352294
rect 439168 352170 439238 352226
rect 439294 352170 439362 352226
rect 439418 352170 439488 352226
rect 439168 352102 439488 352170
rect 439168 352046 439238 352102
rect 439294 352046 439362 352102
rect 439418 352046 439488 352102
rect 439168 351978 439488 352046
rect 439168 351922 439238 351978
rect 439294 351922 439362 351978
rect 439418 351922 439488 351978
rect 439168 351888 439488 351922
rect 469888 352350 470208 352384
rect 469888 352294 469958 352350
rect 470014 352294 470082 352350
rect 470138 352294 470208 352350
rect 469888 352226 470208 352294
rect 469888 352170 469958 352226
rect 470014 352170 470082 352226
rect 470138 352170 470208 352226
rect 469888 352102 470208 352170
rect 469888 352046 469958 352102
rect 470014 352046 470082 352102
rect 470138 352046 470208 352102
rect 469888 351978 470208 352046
rect 469888 351922 469958 351978
rect 470014 351922 470082 351978
rect 470138 351922 470208 351978
rect 469888 351888 470208 351922
rect 500608 352350 500928 352384
rect 500608 352294 500678 352350
rect 500734 352294 500802 352350
rect 500858 352294 500928 352350
rect 500608 352226 500928 352294
rect 500608 352170 500678 352226
rect 500734 352170 500802 352226
rect 500858 352170 500928 352226
rect 500608 352102 500928 352170
rect 500608 352046 500678 352102
rect 500734 352046 500802 352102
rect 500858 352046 500928 352102
rect 500608 351978 500928 352046
rect 500608 351922 500678 351978
rect 500734 351922 500802 351978
rect 500858 351922 500928 351978
rect 500608 351888 500928 351922
rect 24448 346350 24768 346384
rect 24448 346294 24518 346350
rect 24574 346294 24642 346350
rect 24698 346294 24768 346350
rect 24448 346226 24768 346294
rect 24448 346170 24518 346226
rect 24574 346170 24642 346226
rect 24698 346170 24768 346226
rect 24448 346102 24768 346170
rect 24448 346046 24518 346102
rect 24574 346046 24642 346102
rect 24698 346046 24768 346102
rect 24448 345978 24768 346046
rect 24448 345922 24518 345978
rect 24574 345922 24642 345978
rect 24698 345922 24768 345978
rect 24448 345888 24768 345922
rect 55168 346350 55488 346384
rect 55168 346294 55238 346350
rect 55294 346294 55362 346350
rect 55418 346294 55488 346350
rect 55168 346226 55488 346294
rect 55168 346170 55238 346226
rect 55294 346170 55362 346226
rect 55418 346170 55488 346226
rect 55168 346102 55488 346170
rect 55168 346046 55238 346102
rect 55294 346046 55362 346102
rect 55418 346046 55488 346102
rect 55168 345978 55488 346046
rect 55168 345922 55238 345978
rect 55294 345922 55362 345978
rect 55418 345922 55488 345978
rect 55168 345888 55488 345922
rect 85888 346350 86208 346384
rect 85888 346294 85958 346350
rect 86014 346294 86082 346350
rect 86138 346294 86208 346350
rect 85888 346226 86208 346294
rect 85888 346170 85958 346226
rect 86014 346170 86082 346226
rect 86138 346170 86208 346226
rect 85888 346102 86208 346170
rect 85888 346046 85958 346102
rect 86014 346046 86082 346102
rect 86138 346046 86208 346102
rect 85888 345978 86208 346046
rect 85888 345922 85958 345978
rect 86014 345922 86082 345978
rect 86138 345922 86208 345978
rect 85888 345888 86208 345922
rect 116608 346350 116928 346384
rect 116608 346294 116678 346350
rect 116734 346294 116802 346350
rect 116858 346294 116928 346350
rect 116608 346226 116928 346294
rect 116608 346170 116678 346226
rect 116734 346170 116802 346226
rect 116858 346170 116928 346226
rect 116608 346102 116928 346170
rect 116608 346046 116678 346102
rect 116734 346046 116802 346102
rect 116858 346046 116928 346102
rect 116608 345978 116928 346046
rect 116608 345922 116678 345978
rect 116734 345922 116802 345978
rect 116858 345922 116928 345978
rect 116608 345888 116928 345922
rect 147328 346350 147648 346384
rect 147328 346294 147398 346350
rect 147454 346294 147522 346350
rect 147578 346294 147648 346350
rect 147328 346226 147648 346294
rect 147328 346170 147398 346226
rect 147454 346170 147522 346226
rect 147578 346170 147648 346226
rect 147328 346102 147648 346170
rect 147328 346046 147398 346102
rect 147454 346046 147522 346102
rect 147578 346046 147648 346102
rect 147328 345978 147648 346046
rect 147328 345922 147398 345978
rect 147454 345922 147522 345978
rect 147578 345922 147648 345978
rect 147328 345888 147648 345922
rect 178048 346350 178368 346384
rect 178048 346294 178118 346350
rect 178174 346294 178242 346350
rect 178298 346294 178368 346350
rect 178048 346226 178368 346294
rect 178048 346170 178118 346226
rect 178174 346170 178242 346226
rect 178298 346170 178368 346226
rect 178048 346102 178368 346170
rect 178048 346046 178118 346102
rect 178174 346046 178242 346102
rect 178298 346046 178368 346102
rect 178048 345978 178368 346046
rect 178048 345922 178118 345978
rect 178174 345922 178242 345978
rect 178298 345922 178368 345978
rect 178048 345888 178368 345922
rect 208768 346350 209088 346384
rect 208768 346294 208838 346350
rect 208894 346294 208962 346350
rect 209018 346294 209088 346350
rect 208768 346226 209088 346294
rect 208768 346170 208838 346226
rect 208894 346170 208962 346226
rect 209018 346170 209088 346226
rect 208768 346102 209088 346170
rect 208768 346046 208838 346102
rect 208894 346046 208962 346102
rect 209018 346046 209088 346102
rect 208768 345978 209088 346046
rect 208768 345922 208838 345978
rect 208894 345922 208962 345978
rect 209018 345922 209088 345978
rect 208768 345888 209088 345922
rect 239488 346350 239808 346384
rect 239488 346294 239558 346350
rect 239614 346294 239682 346350
rect 239738 346294 239808 346350
rect 239488 346226 239808 346294
rect 239488 346170 239558 346226
rect 239614 346170 239682 346226
rect 239738 346170 239808 346226
rect 239488 346102 239808 346170
rect 239488 346046 239558 346102
rect 239614 346046 239682 346102
rect 239738 346046 239808 346102
rect 239488 345978 239808 346046
rect 239488 345922 239558 345978
rect 239614 345922 239682 345978
rect 239738 345922 239808 345978
rect 239488 345888 239808 345922
rect 270208 346350 270528 346384
rect 270208 346294 270278 346350
rect 270334 346294 270402 346350
rect 270458 346294 270528 346350
rect 270208 346226 270528 346294
rect 270208 346170 270278 346226
rect 270334 346170 270402 346226
rect 270458 346170 270528 346226
rect 270208 346102 270528 346170
rect 270208 346046 270278 346102
rect 270334 346046 270402 346102
rect 270458 346046 270528 346102
rect 270208 345978 270528 346046
rect 270208 345922 270278 345978
rect 270334 345922 270402 345978
rect 270458 345922 270528 345978
rect 270208 345888 270528 345922
rect 300928 346350 301248 346384
rect 300928 346294 300998 346350
rect 301054 346294 301122 346350
rect 301178 346294 301248 346350
rect 300928 346226 301248 346294
rect 300928 346170 300998 346226
rect 301054 346170 301122 346226
rect 301178 346170 301248 346226
rect 300928 346102 301248 346170
rect 300928 346046 300998 346102
rect 301054 346046 301122 346102
rect 301178 346046 301248 346102
rect 300928 345978 301248 346046
rect 300928 345922 300998 345978
rect 301054 345922 301122 345978
rect 301178 345922 301248 345978
rect 300928 345888 301248 345922
rect 331648 346350 331968 346384
rect 331648 346294 331718 346350
rect 331774 346294 331842 346350
rect 331898 346294 331968 346350
rect 331648 346226 331968 346294
rect 331648 346170 331718 346226
rect 331774 346170 331842 346226
rect 331898 346170 331968 346226
rect 331648 346102 331968 346170
rect 331648 346046 331718 346102
rect 331774 346046 331842 346102
rect 331898 346046 331968 346102
rect 331648 345978 331968 346046
rect 331648 345922 331718 345978
rect 331774 345922 331842 345978
rect 331898 345922 331968 345978
rect 331648 345888 331968 345922
rect 362368 346350 362688 346384
rect 362368 346294 362438 346350
rect 362494 346294 362562 346350
rect 362618 346294 362688 346350
rect 362368 346226 362688 346294
rect 362368 346170 362438 346226
rect 362494 346170 362562 346226
rect 362618 346170 362688 346226
rect 362368 346102 362688 346170
rect 362368 346046 362438 346102
rect 362494 346046 362562 346102
rect 362618 346046 362688 346102
rect 362368 345978 362688 346046
rect 362368 345922 362438 345978
rect 362494 345922 362562 345978
rect 362618 345922 362688 345978
rect 362368 345888 362688 345922
rect 393088 346350 393408 346384
rect 393088 346294 393158 346350
rect 393214 346294 393282 346350
rect 393338 346294 393408 346350
rect 393088 346226 393408 346294
rect 393088 346170 393158 346226
rect 393214 346170 393282 346226
rect 393338 346170 393408 346226
rect 393088 346102 393408 346170
rect 393088 346046 393158 346102
rect 393214 346046 393282 346102
rect 393338 346046 393408 346102
rect 393088 345978 393408 346046
rect 393088 345922 393158 345978
rect 393214 345922 393282 345978
rect 393338 345922 393408 345978
rect 393088 345888 393408 345922
rect 423808 346350 424128 346384
rect 423808 346294 423878 346350
rect 423934 346294 424002 346350
rect 424058 346294 424128 346350
rect 423808 346226 424128 346294
rect 423808 346170 423878 346226
rect 423934 346170 424002 346226
rect 424058 346170 424128 346226
rect 423808 346102 424128 346170
rect 423808 346046 423878 346102
rect 423934 346046 424002 346102
rect 424058 346046 424128 346102
rect 423808 345978 424128 346046
rect 423808 345922 423878 345978
rect 423934 345922 424002 345978
rect 424058 345922 424128 345978
rect 423808 345888 424128 345922
rect 454528 346350 454848 346384
rect 454528 346294 454598 346350
rect 454654 346294 454722 346350
rect 454778 346294 454848 346350
rect 454528 346226 454848 346294
rect 454528 346170 454598 346226
rect 454654 346170 454722 346226
rect 454778 346170 454848 346226
rect 454528 346102 454848 346170
rect 454528 346046 454598 346102
rect 454654 346046 454722 346102
rect 454778 346046 454848 346102
rect 454528 345978 454848 346046
rect 454528 345922 454598 345978
rect 454654 345922 454722 345978
rect 454778 345922 454848 345978
rect 454528 345888 454848 345922
rect 485248 346350 485568 346384
rect 485248 346294 485318 346350
rect 485374 346294 485442 346350
rect 485498 346294 485568 346350
rect 485248 346226 485568 346294
rect 485248 346170 485318 346226
rect 485374 346170 485442 346226
rect 485498 346170 485568 346226
rect 485248 346102 485568 346170
rect 485248 346046 485318 346102
rect 485374 346046 485442 346102
rect 485498 346046 485568 346102
rect 485248 345978 485568 346046
rect 485248 345922 485318 345978
rect 485374 345922 485442 345978
rect 485498 345922 485568 345978
rect 485248 345888 485568 345922
rect 515968 346350 516288 346384
rect 515968 346294 516038 346350
rect 516094 346294 516162 346350
rect 516218 346294 516288 346350
rect 515968 346226 516288 346294
rect 515968 346170 516038 346226
rect 516094 346170 516162 346226
rect 516218 346170 516288 346226
rect 515968 346102 516288 346170
rect 515968 346046 516038 346102
rect 516094 346046 516162 346102
rect 516218 346046 516288 346102
rect 515968 345978 516288 346046
rect 515968 345922 516038 345978
rect 516094 345922 516162 345978
rect 516218 345922 516288 345978
rect 515968 345888 516288 345922
rect 525154 346350 525774 363922
rect 525154 346294 525250 346350
rect 525306 346294 525374 346350
rect 525430 346294 525498 346350
rect 525554 346294 525622 346350
rect 525678 346294 525774 346350
rect 525154 346226 525774 346294
rect 525154 346170 525250 346226
rect 525306 346170 525374 346226
rect 525430 346170 525498 346226
rect 525554 346170 525622 346226
rect 525678 346170 525774 346226
rect 525154 346102 525774 346170
rect 525154 346046 525250 346102
rect 525306 346046 525374 346102
rect 525430 346046 525498 346102
rect 525554 346046 525622 346102
rect 525678 346046 525774 346102
rect 525154 345978 525774 346046
rect 525154 345922 525250 345978
rect 525306 345922 525374 345978
rect 525430 345922 525498 345978
rect 525554 345922 525622 345978
rect 525678 345922 525774 345978
rect 6874 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 7494 334350
rect 6874 334226 7494 334294
rect 6874 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 7494 334226
rect 6874 334102 7494 334170
rect 6874 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 7494 334102
rect 6874 333978 7494 334046
rect 6874 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 7494 333978
rect 6874 316350 7494 333922
rect 39808 334350 40128 334384
rect 39808 334294 39878 334350
rect 39934 334294 40002 334350
rect 40058 334294 40128 334350
rect 39808 334226 40128 334294
rect 39808 334170 39878 334226
rect 39934 334170 40002 334226
rect 40058 334170 40128 334226
rect 39808 334102 40128 334170
rect 39808 334046 39878 334102
rect 39934 334046 40002 334102
rect 40058 334046 40128 334102
rect 39808 333978 40128 334046
rect 39808 333922 39878 333978
rect 39934 333922 40002 333978
rect 40058 333922 40128 333978
rect 39808 333888 40128 333922
rect 70528 334350 70848 334384
rect 70528 334294 70598 334350
rect 70654 334294 70722 334350
rect 70778 334294 70848 334350
rect 70528 334226 70848 334294
rect 70528 334170 70598 334226
rect 70654 334170 70722 334226
rect 70778 334170 70848 334226
rect 70528 334102 70848 334170
rect 70528 334046 70598 334102
rect 70654 334046 70722 334102
rect 70778 334046 70848 334102
rect 70528 333978 70848 334046
rect 70528 333922 70598 333978
rect 70654 333922 70722 333978
rect 70778 333922 70848 333978
rect 70528 333888 70848 333922
rect 101248 334350 101568 334384
rect 101248 334294 101318 334350
rect 101374 334294 101442 334350
rect 101498 334294 101568 334350
rect 101248 334226 101568 334294
rect 101248 334170 101318 334226
rect 101374 334170 101442 334226
rect 101498 334170 101568 334226
rect 101248 334102 101568 334170
rect 101248 334046 101318 334102
rect 101374 334046 101442 334102
rect 101498 334046 101568 334102
rect 101248 333978 101568 334046
rect 101248 333922 101318 333978
rect 101374 333922 101442 333978
rect 101498 333922 101568 333978
rect 101248 333888 101568 333922
rect 131968 334350 132288 334384
rect 131968 334294 132038 334350
rect 132094 334294 132162 334350
rect 132218 334294 132288 334350
rect 131968 334226 132288 334294
rect 131968 334170 132038 334226
rect 132094 334170 132162 334226
rect 132218 334170 132288 334226
rect 131968 334102 132288 334170
rect 131968 334046 132038 334102
rect 132094 334046 132162 334102
rect 132218 334046 132288 334102
rect 131968 333978 132288 334046
rect 131968 333922 132038 333978
rect 132094 333922 132162 333978
rect 132218 333922 132288 333978
rect 131968 333888 132288 333922
rect 162688 334350 163008 334384
rect 162688 334294 162758 334350
rect 162814 334294 162882 334350
rect 162938 334294 163008 334350
rect 162688 334226 163008 334294
rect 162688 334170 162758 334226
rect 162814 334170 162882 334226
rect 162938 334170 163008 334226
rect 162688 334102 163008 334170
rect 162688 334046 162758 334102
rect 162814 334046 162882 334102
rect 162938 334046 163008 334102
rect 162688 333978 163008 334046
rect 162688 333922 162758 333978
rect 162814 333922 162882 333978
rect 162938 333922 163008 333978
rect 162688 333888 163008 333922
rect 193408 334350 193728 334384
rect 193408 334294 193478 334350
rect 193534 334294 193602 334350
rect 193658 334294 193728 334350
rect 193408 334226 193728 334294
rect 193408 334170 193478 334226
rect 193534 334170 193602 334226
rect 193658 334170 193728 334226
rect 193408 334102 193728 334170
rect 193408 334046 193478 334102
rect 193534 334046 193602 334102
rect 193658 334046 193728 334102
rect 193408 333978 193728 334046
rect 193408 333922 193478 333978
rect 193534 333922 193602 333978
rect 193658 333922 193728 333978
rect 193408 333888 193728 333922
rect 224128 334350 224448 334384
rect 224128 334294 224198 334350
rect 224254 334294 224322 334350
rect 224378 334294 224448 334350
rect 224128 334226 224448 334294
rect 224128 334170 224198 334226
rect 224254 334170 224322 334226
rect 224378 334170 224448 334226
rect 224128 334102 224448 334170
rect 224128 334046 224198 334102
rect 224254 334046 224322 334102
rect 224378 334046 224448 334102
rect 224128 333978 224448 334046
rect 224128 333922 224198 333978
rect 224254 333922 224322 333978
rect 224378 333922 224448 333978
rect 224128 333888 224448 333922
rect 254848 334350 255168 334384
rect 254848 334294 254918 334350
rect 254974 334294 255042 334350
rect 255098 334294 255168 334350
rect 254848 334226 255168 334294
rect 254848 334170 254918 334226
rect 254974 334170 255042 334226
rect 255098 334170 255168 334226
rect 254848 334102 255168 334170
rect 254848 334046 254918 334102
rect 254974 334046 255042 334102
rect 255098 334046 255168 334102
rect 254848 333978 255168 334046
rect 254848 333922 254918 333978
rect 254974 333922 255042 333978
rect 255098 333922 255168 333978
rect 254848 333888 255168 333922
rect 285568 334350 285888 334384
rect 285568 334294 285638 334350
rect 285694 334294 285762 334350
rect 285818 334294 285888 334350
rect 285568 334226 285888 334294
rect 285568 334170 285638 334226
rect 285694 334170 285762 334226
rect 285818 334170 285888 334226
rect 285568 334102 285888 334170
rect 285568 334046 285638 334102
rect 285694 334046 285762 334102
rect 285818 334046 285888 334102
rect 285568 333978 285888 334046
rect 285568 333922 285638 333978
rect 285694 333922 285762 333978
rect 285818 333922 285888 333978
rect 285568 333888 285888 333922
rect 316288 334350 316608 334384
rect 316288 334294 316358 334350
rect 316414 334294 316482 334350
rect 316538 334294 316608 334350
rect 316288 334226 316608 334294
rect 316288 334170 316358 334226
rect 316414 334170 316482 334226
rect 316538 334170 316608 334226
rect 316288 334102 316608 334170
rect 316288 334046 316358 334102
rect 316414 334046 316482 334102
rect 316538 334046 316608 334102
rect 316288 333978 316608 334046
rect 316288 333922 316358 333978
rect 316414 333922 316482 333978
rect 316538 333922 316608 333978
rect 316288 333888 316608 333922
rect 347008 334350 347328 334384
rect 347008 334294 347078 334350
rect 347134 334294 347202 334350
rect 347258 334294 347328 334350
rect 347008 334226 347328 334294
rect 347008 334170 347078 334226
rect 347134 334170 347202 334226
rect 347258 334170 347328 334226
rect 347008 334102 347328 334170
rect 347008 334046 347078 334102
rect 347134 334046 347202 334102
rect 347258 334046 347328 334102
rect 347008 333978 347328 334046
rect 347008 333922 347078 333978
rect 347134 333922 347202 333978
rect 347258 333922 347328 333978
rect 347008 333888 347328 333922
rect 377728 334350 378048 334384
rect 377728 334294 377798 334350
rect 377854 334294 377922 334350
rect 377978 334294 378048 334350
rect 377728 334226 378048 334294
rect 377728 334170 377798 334226
rect 377854 334170 377922 334226
rect 377978 334170 378048 334226
rect 377728 334102 378048 334170
rect 377728 334046 377798 334102
rect 377854 334046 377922 334102
rect 377978 334046 378048 334102
rect 377728 333978 378048 334046
rect 377728 333922 377798 333978
rect 377854 333922 377922 333978
rect 377978 333922 378048 333978
rect 377728 333888 378048 333922
rect 408448 334350 408768 334384
rect 408448 334294 408518 334350
rect 408574 334294 408642 334350
rect 408698 334294 408768 334350
rect 408448 334226 408768 334294
rect 408448 334170 408518 334226
rect 408574 334170 408642 334226
rect 408698 334170 408768 334226
rect 408448 334102 408768 334170
rect 408448 334046 408518 334102
rect 408574 334046 408642 334102
rect 408698 334046 408768 334102
rect 408448 333978 408768 334046
rect 408448 333922 408518 333978
rect 408574 333922 408642 333978
rect 408698 333922 408768 333978
rect 408448 333888 408768 333922
rect 439168 334350 439488 334384
rect 439168 334294 439238 334350
rect 439294 334294 439362 334350
rect 439418 334294 439488 334350
rect 439168 334226 439488 334294
rect 439168 334170 439238 334226
rect 439294 334170 439362 334226
rect 439418 334170 439488 334226
rect 439168 334102 439488 334170
rect 439168 334046 439238 334102
rect 439294 334046 439362 334102
rect 439418 334046 439488 334102
rect 439168 333978 439488 334046
rect 439168 333922 439238 333978
rect 439294 333922 439362 333978
rect 439418 333922 439488 333978
rect 439168 333888 439488 333922
rect 469888 334350 470208 334384
rect 469888 334294 469958 334350
rect 470014 334294 470082 334350
rect 470138 334294 470208 334350
rect 469888 334226 470208 334294
rect 469888 334170 469958 334226
rect 470014 334170 470082 334226
rect 470138 334170 470208 334226
rect 469888 334102 470208 334170
rect 469888 334046 469958 334102
rect 470014 334046 470082 334102
rect 470138 334046 470208 334102
rect 469888 333978 470208 334046
rect 469888 333922 469958 333978
rect 470014 333922 470082 333978
rect 470138 333922 470208 333978
rect 469888 333888 470208 333922
rect 500608 334350 500928 334384
rect 500608 334294 500678 334350
rect 500734 334294 500802 334350
rect 500858 334294 500928 334350
rect 500608 334226 500928 334294
rect 500608 334170 500678 334226
rect 500734 334170 500802 334226
rect 500858 334170 500928 334226
rect 500608 334102 500928 334170
rect 500608 334046 500678 334102
rect 500734 334046 500802 334102
rect 500858 334046 500928 334102
rect 500608 333978 500928 334046
rect 500608 333922 500678 333978
rect 500734 333922 500802 333978
rect 500858 333922 500928 333978
rect 500608 333888 500928 333922
rect 24448 328350 24768 328384
rect 24448 328294 24518 328350
rect 24574 328294 24642 328350
rect 24698 328294 24768 328350
rect 24448 328226 24768 328294
rect 24448 328170 24518 328226
rect 24574 328170 24642 328226
rect 24698 328170 24768 328226
rect 24448 328102 24768 328170
rect 24448 328046 24518 328102
rect 24574 328046 24642 328102
rect 24698 328046 24768 328102
rect 24448 327978 24768 328046
rect 24448 327922 24518 327978
rect 24574 327922 24642 327978
rect 24698 327922 24768 327978
rect 24448 327888 24768 327922
rect 55168 328350 55488 328384
rect 55168 328294 55238 328350
rect 55294 328294 55362 328350
rect 55418 328294 55488 328350
rect 55168 328226 55488 328294
rect 55168 328170 55238 328226
rect 55294 328170 55362 328226
rect 55418 328170 55488 328226
rect 55168 328102 55488 328170
rect 55168 328046 55238 328102
rect 55294 328046 55362 328102
rect 55418 328046 55488 328102
rect 55168 327978 55488 328046
rect 55168 327922 55238 327978
rect 55294 327922 55362 327978
rect 55418 327922 55488 327978
rect 55168 327888 55488 327922
rect 85888 328350 86208 328384
rect 85888 328294 85958 328350
rect 86014 328294 86082 328350
rect 86138 328294 86208 328350
rect 85888 328226 86208 328294
rect 85888 328170 85958 328226
rect 86014 328170 86082 328226
rect 86138 328170 86208 328226
rect 85888 328102 86208 328170
rect 85888 328046 85958 328102
rect 86014 328046 86082 328102
rect 86138 328046 86208 328102
rect 85888 327978 86208 328046
rect 85888 327922 85958 327978
rect 86014 327922 86082 327978
rect 86138 327922 86208 327978
rect 85888 327888 86208 327922
rect 116608 328350 116928 328384
rect 116608 328294 116678 328350
rect 116734 328294 116802 328350
rect 116858 328294 116928 328350
rect 116608 328226 116928 328294
rect 116608 328170 116678 328226
rect 116734 328170 116802 328226
rect 116858 328170 116928 328226
rect 116608 328102 116928 328170
rect 116608 328046 116678 328102
rect 116734 328046 116802 328102
rect 116858 328046 116928 328102
rect 116608 327978 116928 328046
rect 116608 327922 116678 327978
rect 116734 327922 116802 327978
rect 116858 327922 116928 327978
rect 116608 327888 116928 327922
rect 147328 328350 147648 328384
rect 147328 328294 147398 328350
rect 147454 328294 147522 328350
rect 147578 328294 147648 328350
rect 147328 328226 147648 328294
rect 147328 328170 147398 328226
rect 147454 328170 147522 328226
rect 147578 328170 147648 328226
rect 147328 328102 147648 328170
rect 147328 328046 147398 328102
rect 147454 328046 147522 328102
rect 147578 328046 147648 328102
rect 147328 327978 147648 328046
rect 147328 327922 147398 327978
rect 147454 327922 147522 327978
rect 147578 327922 147648 327978
rect 147328 327888 147648 327922
rect 178048 328350 178368 328384
rect 178048 328294 178118 328350
rect 178174 328294 178242 328350
rect 178298 328294 178368 328350
rect 178048 328226 178368 328294
rect 178048 328170 178118 328226
rect 178174 328170 178242 328226
rect 178298 328170 178368 328226
rect 178048 328102 178368 328170
rect 178048 328046 178118 328102
rect 178174 328046 178242 328102
rect 178298 328046 178368 328102
rect 178048 327978 178368 328046
rect 178048 327922 178118 327978
rect 178174 327922 178242 327978
rect 178298 327922 178368 327978
rect 178048 327888 178368 327922
rect 208768 328350 209088 328384
rect 208768 328294 208838 328350
rect 208894 328294 208962 328350
rect 209018 328294 209088 328350
rect 208768 328226 209088 328294
rect 208768 328170 208838 328226
rect 208894 328170 208962 328226
rect 209018 328170 209088 328226
rect 208768 328102 209088 328170
rect 208768 328046 208838 328102
rect 208894 328046 208962 328102
rect 209018 328046 209088 328102
rect 208768 327978 209088 328046
rect 208768 327922 208838 327978
rect 208894 327922 208962 327978
rect 209018 327922 209088 327978
rect 208768 327888 209088 327922
rect 239488 328350 239808 328384
rect 239488 328294 239558 328350
rect 239614 328294 239682 328350
rect 239738 328294 239808 328350
rect 239488 328226 239808 328294
rect 239488 328170 239558 328226
rect 239614 328170 239682 328226
rect 239738 328170 239808 328226
rect 239488 328102 239808 328170
rect 239488 328046 239558 328102
rect 239614 328046 239682 328102
rect 239738 328046 239808 328102
rect 239488 327978 239808 328046
rect 239488 327922 239558 327978
rect 239614 327922 239682 327978
rect 239738 327922 239808 327978
rect 239488 327888 239808 327922
rect 270208 328350 270528 328384
rect 270208 328294 270278 328350
rect 270334 328294 270402 328350
rect 270458 328294 270528 328350
rect 270208 328226 270528 328294
rect 270208 328170 270278 328226
rect 270334 328170 270402 328226
rect 270458 328170 270528 328226
rect 270208 328102 270528 328170
rect 270208 328046 270278 328102
rect 270334 328046 270402 328102
rect 270458 328046 270528 328102
rect 270208 327978 270528 328046
rect 270208 327922 270278 327978
rect 270334 327922 270402 327978
rect 270458 327922 270528 327978
rect 270208 327888 270528 327922
rect 300928 328350 301248 328384
rect 300928 328294 300998 328350
rect 301054 328294 301122 328350
rect 301178 328294 301248 328350
rect 300928 328226 301248 328294
rect 300928 328170 300998 328226
rect 301054 328170 301122 328226
rect 301178 328170 301248 328226
rect 300928 328102 301248 328170
rect 300928 328046 300998 328102
rect 301054 328046 301122 328102
rect 301178 328046 301248 328102
rect 300928 327978 301248 328046
rect 300928 327922 300998 327978
rect 301054 327922 301122 327978
rect 301178 327922 301248 327978
rect 300928 327888 301248 327922
rect 331648 328350 331968 328384
rect 331648 328294 331718 328350
rect 331774 328294 331842 328350
rect 331898 328294 331968 328350
rect 331648 328226 331968 328294
rect 331648 328170 331718 328226
rect 331774 328170 331842 328226
rect 331898 328170 331968 328226
rect 331648 328102 331968 328170
rect 331648 328046 331718 328102
rect 331774 328046 331842 328102
rect 331898 328046 331968 328102
rect 331648 327978 331968 328046
rect 331648 327922 331718 327978
rect 331774 327922 331842 327978
rect 331898 327922 331968 327978
rect 331648 327888 331968 327922
rect 362368 328350 362688 328384
rect 362368 328294 362438 328350
rect 362494 328294 362562 328350
rect 362618 328294 362688 328350
rect 362368 328226 362688 328294
rect 362368 328170 362438 328226
rect 362494 328170 362562 328226
rect 362618 328170 362688 328226
rect 362368 328102 362688 328170
rect 362368 328046 362438 328102
rect 362494 328046 362562 328102
rect 362618 328046 362688 328102
rect 362368 327978 362688 328046
rect 362368 327922 362438 327978
rect 362494 327922 362562 327978
rect 362618 327922 362688 327978
rect 362368 327888 362688 327922
rect 393088 328350 393408 328384
rect 393088 328294 393158 328350
rect 393214 328294 393282 328350
rect 393338 328294 393408 328350
rect 393088 328226 393408 328294
rect 393088 328170 393158 328226
rect 393214 328170 393282 328226
rect 393338 328170 393408 328226
rect 393088 328102 393408 328170
rect 393088 328046 393158 328102
rect 393214 328046 393282 328102
rect 393338 328046 393408 328102
rect 393088 327978 393408 328046
rect 393088 327922 393158 327978
rect 393214 327922 393282 327978
rect 393338 327922 393408 327978
rect 393088 327888 393408 327922
rect 423808 328350 424128 328384
rect 423808 328294 423878 328350
rect 423934 328294 424002 328350
rect 424058 328294 424128 328350
rect 423808 328226 424128 328294
rect 423808 328170 423878 328226
rect 423934 328170 424002 328226
rect 424058 328170 424128 328226
rect 423808 328102 424128 328170
rect 423808 328046 423878 328102
rect 423934 328046 424002 328102
rect 424058 328046 424128 328102
rect 423808 327978 424128 328046
rect 423808 327922 423878 327978
rect 423934 327922 424002 327978
rect 424058 327922 424128 327978
rect 423808 327888 424128 327922
rect 454528 328350 454848 328384
rect 454528 328294 454598 328350
rect 454654 328294 454722 328350
rect 454778 328294 454848 328350
rect 454528 328226 454848 328294
rect 454528 328170 454598 328226
rect 454654 328170 454722 328226
rect 454778 328170 454848 328226
rect 454528 328102 454848 328170
rect 454528 328046 454598 328102
rect 454654 328046 454722 328102
rect 454778 328046 454848 328102
rect 454528 327978 454848 328046
rect 454528 327922 454598 327978
rect 454654 327922 454722 327978
rect 454778 327922 454848 327978
rect 454528 327888 454848 327922
rect 485248 328350 485568 328384
rect 485248 328294 485318 328350
rect 485374 328294 485442 328350
rect 485498 328294 485568 328350
rect 485248 328226 485568 328294
rect 485248 328170 485318 328226
rect 485374 328170 485442 328226
rect 485498 328170 485568 328226
rect 485248 328102 485568 328170
rect 485248 328046 485318 328102
rect 485374 328046 485442 328102
rect 485498 328046 485568 328102
rect 485248 327978 485568 328046
rect 485248 327922 485318 327978
rect 485374 327922 485442 327978
rect 485498 327922 485568 327978
rect 485248 327888 485568 327922
rect 515968 328350 516288 328384
rect 515968 328294 516038 328350
rect 516094 328294 516162 328350
rect 516218 328294 516288 328350
rect 515968 328226 516288 328294
rect 515968 328170 516038 328226
rect 516094 328170 516162 328226
rect 516218 328170 516288 328226
rect 515968 328102 516288 328170
rect 515968 328046 516038 328102
rect 516094 328046 516162 328102
rect 516218 328046 516288 328102
rect 515968 327978 516288 328046
rect 515968 327922 516038 327978
rect 516094 327922 516162 327978
rect 516218 327922 516288 327978
rect 515968 327888 516288 327922
rect 525154 328350 525774 345922
rect 525154 328294 525250 328350
rect 525306 328294 525374 328350
rect 525430 328294 525498 328350
rect 525554 328294 525622 328350
rect 525678 328294 525774 328350
rect 525154 328226 525774 328294
rect 525154 328170 525250 328226
rect 525306 328170 525374 328226
rect 525430 328170 525498 328226
rect 525554 328170 525622 328226
rect 525678 328170 525774 328226
rect 525154 328102 525774 328170
rect 525154 328046 525250 328102
rect 525306 328046 525374 328102
rect 525430 328046 525498 328102
rect 525554 328046 525622 328102
rect 525678 328046 525774 328102
rect 525154 327978 525774 328046
rect 525154 327922 525250 327978
rect 525306 327922 525374 327978
rect 525430 327922 525498 327978
rect 525554 327922 525622 327978
rect 525678 327922 525774 327978
rect 6874 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 7494 316350
rect 6874 316226 7494 316294
rect 6874 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 7494 316226
rect 6874 316102 7494 316170
rect 6874 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 7494 316102
rect 6874 315978 7494 316046
rect 6874 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 7494 315978
rect 6874 298350 7494 315922
rect 39808 316350 40128 316384
rect 39808 316294 39878 316350
rect 39934 316294 40002 316350
rect 40058 316294 40128 316350
rect 39808 316226 40128 316294
rect 39808 316170 39878 316226
rect 39934 316170 40002 316226
rect 40058 316170 40128 316226
rect 39808 316102 40128 316170
rect 39808 316046 39878 316102
rect 39934 316046 40002 316102
rect 40058 316046 40128 316102
rect 39808 315978 40128 316046
rect 39808 315922 39878 315978
rect 39934 315922 40002 315978
rect 40058 315922 40128 315978
rect 39808 315888 40128 315922
rect 70528 316350 70848 316384
rect 70528 316294 70598 316350
rect 70654 316294 70722 316350
rect 70778 316294 70848 316350
rect 70528 316226 70848 316294
rect 70528 316170 70598 316226
rect 70654 316170 70722 316226
rect 70778 316170 70848 316226
rect 70528 316102 70848 316170
rect 70528 316046 70598 316102
rect 70654 316046 70722 316102
rect 70778 316046 70848 316102
rect 70528 315978 70848 316046
rect 70528 315922 70598 315978
rect 70654 315922 70722 315978
rect 70778 315922 70848 315978
rect 70528 315888 70848 315922
rect 101248 316350 101568 316384
rect 101248 316294 101318 316350
rect 101374 316294 101442 316350
rect 101498 316294 101568 316350
rect 101248 316226 101568 316294
rect 101248 316170 101318 316226
rect 101374 316170 101442 316226
rect 101498 316170 101568 316226
rect 101248 316102 101568 316170
rect 101248 316046 101318 316102
rect 101374 316046 101442 316102
rect 101498 316046 101568 316102
rect 101248 315978 101568 316046
rect 101248 315922 101318 315978
rect 101374 315922 101442 315978
rect 101498 315922 101568 315978
rect 101248 315888 101568 315922
rect 131968 316350 132288 316384
rect 131968 316294 132038 316350
rect 132094 316294 132162 316350
rect 132218 316294 132288 316350
rect 131968 316226 132288 316294
rect 131968 316170 132038 316226
rect 132094 316170 132162 316226
rect 132218 316170 132288 316226
rect 131968 316102 132288 316170
rect 131968 316046 132038 316102
rect 132094 316046 132162 316102
rect 132218 316046 132288 316102
rect 131968 315978 132288 316046
rect 131968 315922 132038 315978
rect 132094 315922 132162 315978
rect 132218 315922 132288 315978
rect 131968 315888 132288 315922
rect 162688 316350 163008 316384
rect 162688 316294 162758 316350
rect 162814 316294 162882 316350
rect 162938 316294 163008 316350
rect 162688 316226 163008 316294
rect 162688 316170 162758 316226
rect 162814 316170 162882 316226
rect 162938 316170 163008 316226
rect 162688 316102 163008 316170
rect 162688 316046 162758 316102
rect 162814 316046 162882 316102
rect 162938 316046 163008 316102
rect 162688 315978 163008 316046
rect 162688 315922 162758 315978
rect 162814 315922 162882 315978
rect 162938 315922 163008 315978
rect 162688 315888 163008 315922
rect 193408 316350 193728 316384
rect 193408 316294 193478 316350
rect 193534 316294 193602 316350
rect 193658 316294 193728 316350
rect 193408 316226 193728 316294
rect 193408 316170 193478 316226
rect 193534 316170 193602 316226
rect 193658 316170 193728 316226
rect 193408 316102 193728 316170
rect 193408 316046 193478 316102
rect 193534 316046 193602 316102
rect 193658 316046 193728 316102
rect 193408 315978 193728 316046
rect 193408 315922 193478 315978
rect 193534 315922 193602 315978
rect 193658 315922 193728 315978
rect 193408 315888 193728 315922
rect 224128 316350 224448 316384
rect 224128 316294 224198 316350
rect 224254 316294 224322 316350
rect 224378 316294 224448 316350
rect 224128 316226 224448 316294
rect 224128 316170 224198 316226
rect 224254 316170 224322 316226
rect 224378 316170 224448 316226
rect 224128 316102 224448 316170
rect 224128 316046 224198 316102
rect 224254 316046 224322 316102
rect 224378 316046 224448 316102
rect 224128 315978 224448 316046
rect 224128 315922 224198 315978
rect 224254 315922 224322 315978
rect 224378 315922 224448 315978
rect 224128 315888 224448 315922
rect 254848 316350 255168 316384
rect 254848 316294 254918 316350
rect 254974 316294 255042 316350
rect 255098 316294 255168 316350
rect 254848 316226 255168 316294
rect 254848 316170 254918 316226
rect 254974 316170 255042 316226
rect 255098 316170 255168 316226
rect 254848 316102 255168 316170
rect 254848 316046 254918 316102
rect 254974 316046 255042 316102
rect 255098 316046 255168 316102
rect 254848 315978 255168 316046
rect 254848 315922 254918 315978
rect 254974 315922 255042 315978
rect 255098 315922 255168 315978
rect 254848 315888 255168 315922
rect 285568 316350 285888 316384
rect 285568 316294 285638 316350
rect 285694 316294 285762 316350
rect 285818 316294 285888 316350
rect 285568 316226 285888 316294
rect 285568 316170 285638 316226
rect 285694 316170 285762 316226
rect 285818 316170 285888 316226
rect 285568 316102 285888 316170
rect 285568 316046 285638 316102
rect 285694 316046 285762 316102
rect 285818 316046 285888 316102
rect 285568 315978 285888 316046
rect 285568 315922 285638 315978
rect 285694 315922 285762 315978
rect 285818 315922 285888 315978
rect 285568 315888 285888 315922
rect 316288 316350 316608 316384
rect 316288 316294 316358 316350
rect 316414 316294 316482 316350
rect 316538 316294 316608 316350
rect 316288 316226 316608 316294
rect 316288 316170 316358 316226
rect 316414 316170 316482 316226
rect 316538 316170 316608 316226
rect 316288 316102 316608 316170
rect 316288 316046 316358 316102
rect 316414 316046 316482 316102
rect 316538 316046 316608 316102
rect 316288 315978 316608 316046
rect 316288 315922 316358 315978
rect 316414 315922 316482 315978
rect 316538 315922 316608 315978
rect 316288 315888 316608 315922
rect 347008 316350 347328 316384
rect 347008 316294 347078 316350
rect 347134 316294 347202 316350
rect 347258 316294 347328 316350
rect 347008 316226 347328 316294
rect 347008 316170 347078 316226
rect 347134 316170 347202 316226
rect 347258 316170 347328 316226
rect 347008 316102 347328 316170
rect 347008 316046 347078 316102
rect 347134 316046 347202 316102
rect 347258 316046 347328 316102
rect 347008 315978 347328 316046
rect 347008 315922 347078 315978
rect 347134 315922 347202 315978
rect 347258 315922 347328 315978
rect 347008 315888 347328 315922
rect 377728 316350 378048 316384
rect 377728 316294 377798 316350
rect 377854 316294 377922 316350
rect 377978 316294 378048 316350
rect 377728 316226 378048 316294
rect 377728 316170 377798 316226
rect 377854 316170 377922 316226
rect 377978 316170 378048 316226
rect 377728 316102 378048 316170
rect 377728 316046 377798 316102
rect 377854 316046 377922 316102
rect 377978 316046 378048 316102
rect 377728 315978 378048 316046
rect 377728 315922 377798 315978
rect 377854 315922 377922 315978
rect 377978 315922 378048 315978
rect 377728 315888 378048 315922
rect 408448 316350 408768 316384
rect 408448 316294 408518 316350
rect 408574 316294 408642 316350
rect 408698 316294 408768 316350
rect 408448 316226 408768 316294
rect 408448 316170 408518 316226
rect 408574 316170 408642 316226
rect 408698 316170 408768 316226
rect 408448 316102 408768 316170
rect 408448 316046 408518 316102
rect 408574 316046 408642 316102
rect 408698 316046 408768 316102
rect 408448 315978 408768 316046
rect 408448 315922 408518 315978
rect 408574 315922 408642 315978
rect 408698 315922 408768 315978
rect 408448 315888 408768 315922
rect 439168 316350 439488 316384
rect 439168 316294 439238 316350
rect 439294 316294 439362 316350
rect 439418 316294 439488 316350
rect 439168 316226 439488 316294
rect 439168 316170 439238 316226
rect 439294 316170 439362 316226
rect 439418 316170 439488 316226
rect 439168 316102 439488 316170
rect 439168 316046 439238 316102
rect 439294 316046 439362 316102
rect 439418 316046 439488 316102
rect 439168 315978 439488 316046
rect 439168 315922 439238 315978
rect 439294 315922 439362 315978
rect 439418 315922 439488 315978
rect 439168 315888 439488 315922
rect 469888 316350 470208 316384
rect 469888 316294 469958 316350
rect 470014 316294 470082 316350
rect 470138 316294 470208 316350
rect 469888 316226 470208 316294
rect 469888 316170 469958 316226
rect 470014 316170 470082 316226
rect 470138 316170 470208 316226
rect 469888 316102 470208 316170
rect 469888 316046 469958 316102
rect 470014 316046 470082 316102
rect 470138 316046 470208 316102
rect 469888 315978 470208 316046
rect 469888 315922 469958 315978
rect 470014 315922 470082 315978
rect 470138 315922 470208 315978
rect 469888 315888 470208 315922
rect 500608 316350 500928 316384
rect 500608 316294 500678 316350
rect 500734 316294 500802 316350
rect 500858 316294 500928 316350
rect 500608 316226 500928 316294
rect 500608 316170 500678 316226
rect 500734 316170 500802 316226
rect 500858 316170 500928 316226
rect 500608 316102 500928 316170
rect 500608 316046 500678 316102
rect 500734 316046 500802 316102
rect 500858 316046 500928 316102
rect 500608 315978 500928 316046
rect 500608 315922 500678 315978
rect 500734 315922 500802 315978
rect 500858 315922 500928 315978
rect 500608 315888 500928 315922
rect 24448 310350 24768 310384
rect 24448 310294 24518 310350
rect 24574 310294 24642 310350
rect 24698 310294 24768 310350
rect 24448 310226 24768 310294
rect 24448 310170 24518 310226
rect 24574 310170 24642 310226
rect 24698 310170 24768 310226
rect 24448 310102 24768 310170
rect 24448 310046 24518 310102
rect 24574 310046 24642 310102
rect 24698 310046 24768 310102
rect 24448 309978 24768 310046
rect 24448 309922 24518 309978
rect 24574 309922 24642 309978
rect 24698 309922 24768 309978
rect 24448 309888 24768 309922
rect 55168 310350 55488 310384
rect 55168 310294 55238 310350
rect 55294 310294 55362 310350
rect 55418 310294 55488 310350
rect 55168 310226 55488 310294
rect 55168 310170 55238 310226
rect 55294 310170 55362 310226
rect 55418 310170 55488 310226
rect 55168 310102 55488 310170
rect 55168 310046 55238 310102
rect 55294 310046 55362 310102
rect 55418 310046 55488 310102
rect 55168 309978 55488 310046
rect 55168 309922 55238 309978
rect 55294 309922 55362 309978
rect 55418 309922 55488 309978
rect 55168 309888 55488 309922
rect 85888 310350 86208 310384
rect 85888 310294 85958 310350
rect 86014 310294 86082 310350
rect 86138 310294 86208 310350
rect 85888 310226 86208 310294
rect 85888 310170 85958 310226
rect 86014 310170 86082 310226
rect 86138 310170 86208 310226
rect 85888 310102 86208 310170
rect 85888 310046 85958 310102
rect 86014 310046 86082 310102
rect 86138 310046 86208 310102
rect 85888 309978 86208 310046
rect 85888 309922 85958 309978
rect 86014 309922 86082 309978
rect 86138 309922 86208 309978
rect 85888 309888 86208 309922
rect 116608 310350 116928 310384
rect 116608 310294 116678 310350
rect 116734 310294 116802 310350
rect 116858 310294 116928 310350
rect 116608 310226 116928 310294
rect 116608 310170 116678 310226
rect 116734 310170 116802 310226
rect 116858 310170 116928 310226
rect 116608 310102 116928 310170
rect 116608 310046 116678 310102
rect 116734 310046 116802 310102
rect 116858 310046 116928 310102
rect 116608 309978 116928 310046
rect 116608 309922 116678 309978
rect 116734 309922 116802 309978
rect 116858 309922 116928 309978
rect 116608 309888 116928 309922
rect 147328 310350 147648 310384
rect 147328 310294 147398 310350
rect 147454 310294 147522 310350
rect 147578 310294 147648 310350
rect 147328 310226 147648 310294
rect 147328 310170 147398 310226
rect 147454 310170 147522 310226
rect 147578 310170 147648 310226
rect 147328 310102 147648 310170
rect 147328 310046 147398 310102
rect 147454 310046 147522 310102
rect 147578 310046 147648 310102
rect 147328 309978 147648 310046
rect 147328 309922 147398 309978
rect 147454 309922 147522 309978
rect 147578 309922 147648 309978
rect 147328 309888 147648 309922
rect 178048 310350 178368 310384
rect 178048 310294 178118 310350
rect 178174 310294 178242 310350
rect 178298 310294 178368 310350
rect 178048 310226 178368 310294
rect 178048 310170 178118 310226
rect 178174 310170 178242 310226
rect 178298 310170 178368 310226
rect 178048 310102 178368 310170
rect 178048 310046 178118 310102
rect 178174 310046 178242 310102
rect 178298 310046 178368 310102
rect 178048 309978 178368 310046
rect 178048 309922 178118 309978
rect 178174 309922 178242 309978
rect 178298 309922 178368 309978
rect 178048 309888 178368 309922
rect 208768 310350 209088 310384
rect 208768 310294 208838 310350
rect 208894 310294 208962 310350
rect 209018 310294 209088 310350
rect 208768 310226 209088 310294
rect 208768 310170 208838 310226
rect 208894 310170 208962 310226
rect 209018 310170 209088 310226
rect 208768 310102 209088 310170
rect 208768 310046 208838 310102
rect 208894 310046 208962 310102
rect 209018 310046 209088 310102
rect 208768 309978 209088 310046
rect 208768 309922 208838 309978
rect 208894 309922 208962 309978
rect 209018 309922 209088 309978
rect 208768 309888 209088 309922
rect 239488 310350 239808 310384
rect 239488 310294 239558 310350
rect 239614 310294 239682 310350
rect 239738 310294 239808 310350
rect 239488 310226 239808 310294
rect 239488 310170 239558 310226
rect 239614 310170 239682 310226
rect 239738 310170 239808 310226
rect 239488 310102 239808 310170
rect 239488 310046 239558 310102
rect 239614 310046 239682 310102
rect 239738 310046 239808 310102
rect 239488 309978 239808 310046
rect 239488 309922 239558 309978
rect 239614 309922 239682 309978
rect 239738 309922 239808 309978
rect 239488 309888 239808 309922
rect 270208 310350 270528 310384
rect 270208 310294 270278 310350
rect 270334 310294 270402 310350
rect 270458 310294 270528 310350
rect 270208 310226 270528 310294
rect 270208 310170 270278 310226
rect 270334 310170 270402 310226
rect 270458 310170 270528 310226
rect 270208 310102 270528 310170
rect 270208 310046 270278 310102
rect 270334 310046 270402 310102
rect 270458 310046 270528 310102
rect 270208 309978 270528 310046
rect 270208 309922 270278 309978
rect 270334 309922 270402 309978
rect 270458 309922 270528 309978
rect 270208 309888 270528 309922
rect 300928 310350 301248 310384
rect 300928 310294 300998 310350
rect 301054 310294 301122 310350
rect 301178 310294 301248 310350
rect 300928 310226 301248 310294
rect 300928 310170 300998 310226
rect 301054 310170 301122 310226
rect 301178 310170 301248 310226
rect 300928 310102 301248 310170
rect 300928 310046 300998 310102
rect 301054 310046 301122 310102
rect 301178 310046 301248 310102
rect 300928 309978 301248 310046
rect 300928 309922 300998 309978
rect 301054 309922 301122 309978
rect 301178 309922 301248 309978
rect 300928 309888 301248 309922
rect 331648 310350 331968 310384
rect 331648 310294 331718 310350
rect 331774 310294 331842 310350
rect 331898 310294 331968 310350
rect 331648 310226 331968 310294
rect 331648 310170 331718 310226
rect 331774 310170 331842 310226
rect 331898 310170 331968 310226
rect 331648 310102 331968 310170
rect 331648 310046 331718 310102
rect 331774 310046 331842 310102
rect 331898 310046 331968 310102
rect 331648 309978 331968 310046
rect 331648 309922 331718 309978
rect 331774 309922 331842 309978
rect 331898 309922 331968 309978
rect 331648 309888 331968 309922
rect 362368 310350 362688 310384
rect 362368 310294 362438 310350
rect 362494 310294 362562 310350
rect 362618 310294 362688 310350
rect 362368 310226 362688 310294
rect 362368 310170 362438 310226
rect 362494 310170 362562 310226
rect 362618 310170 362688 310226
rect 362368 310102 362688 310170
rect 362368 310046 362438 310102
rect 362494 310046 362562 310102
rect 362618 310046 362688 310102
rect 362368 309978 362688 310046
rect 362368 309922 362438 309978
rect 362494 309922 362562 309978
rect 362618 309922 362688 309978
rect 362368 309888 362688 309922
rect 393088 310350 393408 310384
rect 393088 310294 393158 310350
rect 393214 310294 393282 310350
rect 393338 310294 393408 310350
rect 393088 310226 393408 310294
rect 393088 310170 393158 310226
rect 393214 310170 393282 310226
rect 393338 310170 393408 310226
rect 393088 310102 393408 310170
rect 393088 310046 393158 310102
rect 393214 310046 393282 310102
rect 393338 310046 393408 310102
rect 393088 309978 393408 310046
rect 393088 309922 393158 309978
rect 393214 309922 393282 309978
rect 393338 309922 393408 309978
rect 393088 309888 393408 309922
rect 423808 310350 424128 310384
rect 423808 310294 423878 310350
rect 423934 310294 424002 310350
rect 424058 310294 424128 310350
rect 423808 310226 424128 310294
rect 423808 310170 423878 310226
rect 423934 310170 424002 310226
rect 424058 310170 424128 310226
rect 423808 310102 424128 310170
rect 423808 310046 423878 310102
rect 423934 310046 424002 310102
rect 424058 310046 424128 310102
rect 423808 309978 424128 310046
rect 423808 309922 423878 309978
rect 423934 309922 424002 309978
rect 424058 309922 424128 309978
rect 423808 309888 424128 309922
rect 454528 310350 454848 310384
rect 454528 310294 454598 310350
rect 454654 310294 454722 310350
rect 454778 310294 454848 310350
rect 454528 310226 454848 310294
rect 454528 310170 454598 310226
rect 454654 310170 454722 310226
rect 454778 310170 454848 310226
rect 454528 310102 454848 310170
rect 454528 310046 454598 310102
rect 454654 310046 454722 310102
rect 454778 310046 454848 310102
rect 454528 309978 454848 310046
rect 454528 309922 454598 309978
rect 454654 309922 454722 309978
rect 454778 309922 454848 309978
rect 454528 309888 454848 309922
rect 485248 310350 485568 310384
rect 485248 310294 485318 310350
rect 485374 310294 485442 310350
rect 485498 310294 485568 310350
rect 485248 310226 485568 310294
rect 485248 310170 485318 310226
rect 485374 310170 485442 310226
rect 485498 310170 485568 310226
rect 485248 310102 485568 310170
rect 485248 310046 485318 310102
rect 485374 310046 485442 310102
rect 485498 310046 485568 310102
rect 485248 309978 485568 310046
rect 485248 309922 485318 309978
rect 485374 309922 485442 309978
rect 485498 309922 485568 309978
rect 485248 309888 485568 309922
rect 515968 310350 516288 310384
rect 515968 310294 516038 310350
rect 516094 310294 516162 310350
rect 516218 310294 516288 310350
rect 515968 310226 516288 310294
rect 515968 310170 516038 310226
rect 516094 310170 516162 310226
rect 516218 310170 516288 310226
rect 515968 310102 516288 310170
rect 515968 310046 516038 310102
rect 516094 310046 516162 310102
rect 516218 310046 516288 310102
rect 515968 309978 516288 310046
rect 515968 309922 516038 309978
rect 516094 309922 516162 309978
rect 516218 309922 516288 309978
rect 515968 309888 516288 309922
rect 525154 310350 525774 327922
rect 525154 310294 525250 310350
rect 525306 310294 525374 310350
rect 525430 310294 525498 310350
rect 525554 310294 525622 310350
rect 525678 310294 525774 310350
rect 525154 310226 525774 310294
rect 525154 310170 525250 310226
rect 525306 310170 525374 310226
rect 525430 310170 525498 310226
rect 525554 310170 525622 310226
rect 525678 310170 525774 310226
rect 525154 310102 525774 310170
rect 525154 310046 525250 310102
rect 525306 310046 525374 310102
rect 525430 310046 525498 310102
rect 525554 310046 525622 310102
rect 525678 310046 525774 310102
rect 525154 309978 525774 310046
rect 525154 309922 525250 309978
rect 525306 309922 525374 309978
rect 525430 309922 525498 309978
rect 525554 309922 525622 309978
rect 525678 309922 525774 309978
rect 6874 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 7494 298350
rect 6874 298226 7494 298294
rect 6874 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 7494 298226
rect 6874 298102 7494 298170
rect 6874 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 7494 298102
rect 6874 297978 7494 298046
rect 6874 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 7494 297978
rect 6874 280350 7494 297922
rect 39808 298350 40128 298384
rect 39808 298294 39878 298350
rect 39934 298294 40002 298350
rect 40058 298294 40128 298350
rect 39808 298226 40128 298294
rect 39808 298170 39878 298226
rect 39934 298170 40002 298226
rect 40058 298170 40128 298226
rect 39808 298102 40128 298170
rect 39808 298046 39878 298102
rect 39934 298046 40002 298102
rect 40058 298046 40128 298102
rect 39808 297978 40128 298046
rect 39808 297922 39878 297978
rect 39934 297922 40002 297978
rect 40058 297922 40128 297978
rect 39808 297888 40128 297922
rect 70528 298350 70848 298384
rect 70528 298294 70598 298350
rect 70654 298294 70722 298350
rect 70778 298294 70848 298350
rect 70528 298226 70848 298294
rect 70528 298170 70598 298226
rect 70654 298170 70722 298226
rect 70778 298170 70848 298226
rect 70528 298102 70848 298170
rect 70528 298046 70598 298102
rect 70654 298046 70722 298102
rect 70778 298046 70848 298102
rect 70528 297978 70848 298046
rect 70528 297922 70598 297978
rect 70654 297922 70722 297978
rect 70778 297922 70848 297978
rect 70528 297888 70848 297922
rect 101248 298350 101568 298384
rect 101248 298294 101318 298350
rect 101374 298294 101442 298350
rect 101498 298294 101568 298350
rect 101248 298226 101568 298294
rect 101248 298170 101318 298226
rect 101374 298170 101442 298226
rect 101498 298170 101568 298226
rect 101248 298102 101568 298170
rect 101248 298046 101318 298102
rect 101374 298046 101442 298102
rect 101498 298046 101568 298102
rect 101248 297978 101568 298046
rect 101248 297922 101318 297978
rect 101374 297922 101442 297978
rect 101498 297922 101568 297978
rect 101248 297888 101568 297922
rect 131968 298350 132288 298384
rect 131968 298294 132038 298350
rect 132094 298294 132162 298350
rect 132218 298294 132288 298350
rect 131968 298226 132288 298294
rect 131968 298170 132038 298226
rect 132094 298170 132162 298226
rect 132218 298170 132288 298226
rect 131968 298102 132288 298170
rect 131968 298046 132038 298102
rect 132094 298046 132162 298102
rect 132218 298046 132288 298102
rect 131968 297978 132288 298046
rect 131968 297922 132038 297978
rect 132094 297922 132162 297978
rect 132218 297922 132288 297978
rect 131968 297888 132288 297922
rect 162688 298350 163008 298384
rect 162688 298294 162758 298350
rect 162814 298294 162882 298350
rect 162938 298294 163008 298350
rect 162688 298226 163008 298294
rect 162688 298170 162758 298226
rect 162814 298170 162882 298226
rect 162938 298170 163008 298226
rect 162688 298102 163008 298170
rect 162688 298046 162758 298102
rect 162814 298046 162882 298102
rect 162938 298046 163008 298102
rect 162688 297978 163008 298046
rect 162688 297922 162758 297978
rect 162814 297922 162882 297978
rect 162938 297922 163008 297978
rect 162688 297888 163008 297922
rect 193408 298350 193728 298384
rect 193408 298294 193478 298350
rect 193534 298294 193602 298350
rect 193658 298294 193728 298350
rect 193408 298226 193728 298294
rect 193408 298170 193478 298226
rect 193534 298170 193602 298226
rect 193658 298170 193728 298226
rect 193408 298102 193728 298170
rect 193408 298046 193478 298102
rect 193534 298046 193602 298102
rect 193658 298046 193728 298102
rect 193408 297978 193728 298046
rect 193408 297922 193478 297978
rect 193534 297922 193602 297978
rect 193658 297922 193728 297978
rect 193408 297888 193728 297922
rect 224128 298350 224448 298384
rect 224128 298294 224198 298350
rect 224254 298294 224322 298350
rect 224378 298294 224448 298350
rect 224128 298226 224448 298294
rect 224128 298170 224198 298226
rect 224254 298170 224322 298226
rect 224378 298170 224448 298226
rect 224128 298102 224448 298170
rect 224128 298046 224198 298102
rect 224254 298046 224322 298102
rect 224378 298046 224448 298102
rect 224128 297978 224448 298046
rect 224128 297922 224198 297978
rect 224254 297922 224322 297978
rect 224378 297922 224448 297978
rect 224128 297888 224448 297922
rect 254848 298350 255168 298384
rect 254848 298294 254918 298350
rect 254974 298294 255042 298350
rect 255098 298294 255168 298350
rect 254848 298226 255168 298294
rect 254848 298170 254918 298226
rect 254974 298170 255042 298226
rect 255098 298170 255168 298226
rect 254848 298102 255168 298170
rect 254848 298046 254918 298102
rect 254974 298046 255042 298102
rect 255098 298046 255168 298102
rect 254848 297978 255168 298046
rect 254848 297922 254918 297978
rect 254974 297922 255042 297978
rect 255098 297922 255168 297978
rect 254848 297888 255168 297922
rect 285568 298350 285888 298384
rect 285568 298294 285638 298350
rect 285694 298294 285762 298350
rect 285818 298294 285888 298350
rect 285568 298226 285888 298294
rect 285568 298170 285638 298226
rect 285694 298170 285762 298226
rect 285818 298170 285888 298226
rect 285568 298102 285888 298170
rect 285568 298046 285638 298102
rect 285694 298046 285762 298102
rect 285818 298046 285888 298102
rect 285568 297978 285888 298046
rect 285568 297922 285638 297978
rect 285694 297922 285762 297978
rect 285818 297922 285888 297978
rect 285568 297888 285888 297922
rect 316288 298350 316608 298384
rect 316288 298294 316358 298350
rect 316414 298294 316482 298350
rect 316538 298294 316608 298350
rect 316288 298226 316608 298294
rect 316288 298170 316358 298226
rect 316414 298170 316482 298226
rect 316538 298170 316608 298226
rect 316288 298102 316608 298170
rect 316288 298046 316358 298102
rect 316414 298046 316482 298102
rect 316538 298046 316608 298102
rect 316288 297978 316608 298046
rect 316288 297922 316358 297978
rect 316414 297922 316482 297978
rect 316538 297922 316608 297978
rect 316288 297888 316608 297922
rect 347008 298350 347328 298384
rect 347008 298294 347078 298350
rect 347134 298294 347202 298350
rect 347258 298294 347328 298350
rect 347008 298226 347328 298294
rect 347008 298170 347078 298226
rect 347134 298170 347202 298226
rect 347258 298170 347328 298226
rect 347008 298102 347328 298170
rect 347008 298046 347078 298102
rect 347134 298046 347202 298102
rect 347258 298046 347328 298102
rect 347008 297978 347328 298046
rect 347008 297922 347078 297978
rect 347134 297922 347202 297978
rect 347258 297922 347328 297978
rect 347008 297888 347328 297922
rect 377728 298350 378048 298384
rect 377728 298294 377798 298350
rect 377854 298294 377922 298350
rect 377978 298294 378048 298350
rect 377728 298226 378048 298294
rect 377728 298170 377798 298226
rect 377854 298170 377922 298226
rect 377978 298170 378048 298226
rect 377728 298102 378048 298170
rect 377728 298046 377798 298102
rect 377854 298046 377922 298102
rect 377978 298046 378048 298102
rect 377728 297978 378048 298046
rect 377728 297922 377798 297978
rect 377854 297922 377922 297978
rect 377978 297922 378048 297978
rect 377728 297888 378048 297922
rect 408448 298350 408768 298384
rect 408448 298294 408518 298350
rect 408574 298294 408642 298350
rect 408698 298294 408768 298350
rect 408448 298226 408768 298294
rect 408448 298170 408518 298226
rect 408574 298170 408642 298226
rect 408698 298170 408768 298226
rect 408448 298102 408768 298170
rect 408448 298046 408518 298102
rect 408574 298046 408642 298102
rect 408698 298046 408768 298102
rect 408448 297978 408768 298046
rect 408448 297922 408518 297978
rect 408574 297922 408642 297978
rect 408698 297922 408768 297978
rect 408448 297888 408768 297922
rect 439168 298350 439488 298384
rect 439168 298294 439238 298350
rect 439294 298294 439362 298350
rect 439418 298294 439488 298350
rect 439168 298226 439488 298294
rect 439168 298170 439238 298226
rect 439294 298170 439362 298226
rect 439418 298170 439488 298226
rect 439168 298102 439488 298170
rect 439168 298046 439238 298102
rect 439294 298046 439362 298102
rect 439418 298046 439488 298102
rect 439168 297978 439488 298046
rect 439168 297922 439238 297978
rect 439294 297922 439362 297978
rect 439418 297922 439488 297978
rect 439168 297888 439488 297922
rect 469888 298350 470208 298384
rect 469888 298294 469958 298350
rect 470014 298294 470082 298350
rect 470138 298294 470208 298350
rect 469888 298226 470208 298294
rect 469888 298170 469958 298226
rect 470014 298170 470082 298226
rect 470138 298170 470208 298226
rect 469888 298102 470208 298170
rect 469888 298046 469958 298102
rect 470014 298046 470082 298102
rect 470138 298046 470208 298102
rect 469888 297978 470208 298046
rect 469888 297922 469958 297978
rect 470014 297922 470082 297978
rect 470138 297922 470208 297978
rect 469888 297888 470208 297922
rect 500608 298350 500928 298384
rect 500608 298294 500678 298350
rect 500734 298294 500802 298350
rect 500858 298294 500928 298350
rect 500608 298226 500928 298294
rect 500608 298170 500678 298226
rect 500734 298170 500802 298226
rect 500858 298170 500928 298226
rect 500608 298102 500928 298170
rect 500608 298046 500678 298102
rect 500734 298046 500802 298102
rect 500858 298046 500928 298102
rect 500608 297978 500928 298046
rect 500608 297922 500678 297978
rect 500734 297922 500802 297978
rect 500858 297922 500928 297978
rect 500608 297888 500928 297922
rect 24448 292350 24768 292384
rect 24448 292294 24518 292350
rect 24574 292294 24642 292350
rect 24698 292294 24768 292350
rect 24448 292226 24768 292294
rect 24448 292170 24518 292226
rect 24574 292170 24642 292226
rect 24698 292170 24768 292226
rect 24448 292102 24768 292170
rect 24448 292046 24518 292102
rect 24574 292046 24642 292102
rect 24698 292046 24768 292102
rect 24448 291978 24768 292046
rect 24448 291922 24518 291978
rect 24574 291922 24642 291978
rect 24698 291922 24768 291978
rect 24448 291888 24768 291922
rect 55168 292350 55488 292384
rect 55168 292294 55238 292350
rect 55294 292294 55362 292350
rect 55418 292294 55488 292350
rect 55168 292226 55488 292294
rect 55168 292170 55238 292226
rect 55294 292170 55362 292226
rect 55418 292170 55488 292226
rect 55168 292102 55488 292170
rect 55168 292046 55238 292102
rect 55294 292046 55362 292102
rect 55418 292046 55488 292102
rect 55168 291978 55488 292046
rect 55168 291922 55238 291978
rect 55294 291922 55362 291978
rect 55418 291922 55488 291978
rect 55168 291888 55488 291922
rect 85888 292350 86208 292384
rect 85888 292294 85958 292350
rect 86014 292294 86082 292350
rect 86138 292294 86208 292350
rect 85888 292226 86208 292294
rect 85888 292170 85958 292226
rect 86014 292170 86082 292226
rect 86138 292170 86208 292226
rect 85888 292102 86208 292170
rect 85888 292046 85958 292102
rect 86014 292046 86082 292102
rect 86138 292046 86208 292102
rect 85888 291978 86208 292046
rect 85888 291922 85958 291978
rect 86014 291922 86082 291978
rect 86138 291922 86208 291978
rect 85888 291888 86208 291922
rect 116608 292350 116928 292384
rect 116608 292294 116678 292350
rect 116734 292294 116802 292350
rect 116858 292294 116928 292350
rect 116608 292226 116928 292294
rect 116608 292170 116678 292226
rect 116734 292170 116802 292226
rect 116858 292170 116928 292226
rect 116608 292102 116928 292170
rect 116608 292046 116678 292102
rect 116734 292046 116802 292102
rect 116858 292046 116928 292102
rect 116608 291978 116928 292046
rect 116608 291922 116678 291978
rect 116734 291922 116802 291978
rect 116858 291922 116928 291978
rect 116608 291888 116928 291922
rect 147328 292350 147648 292384
rect 147328 292294 147398 292350
rect 147454 292294 147522 292350
rect 147578 292294 147648 292350
rect 147328 292226 147648 292294
rect 147328 292170 147398 292226
rect 147454 292170 147522 292226
rect 147578 292170 147648 292226
rect 147328 292102 147648 292170
rect 147328 292046 147398 292102
rect 147454 292046 147522 292102
rect 147578 292046 147648 292102
rect 147328 291978 147648 292046
rect 147328 291922 147398 291978
rect 147454 291922 147522 291978
rect 147578 291922 147648 291978
rect 147328 291888 147648 291922
rect 178048 292350 178368 292384
rect 178048 292294 178118 292350
rect 178174 292294 178242 292350
rect 178298 292294 178368 292350
rect 178048 292226 178368 292294
rect 178048 292170 178118 292226
rect 178174 292170 178242 292226
rect 178298 292170 178368 292226
rect 178048 292102 178368 292170
rect 178048 292046 178118 292102
rect 178174 292046 178242 292102
rect 178298 292046 178368 292102
rect 178048 291978 178368 292046
rect 178048 291922 178118 291978
rect 178174 291922 178242 291978
rect 178298 291922 178368 291978
rect 178048 291888 178368 291922
rect 208768 292350 209088 292384
rect 208768 292294 208838 292350
rect 208894 292294 208962 292350
rect 209018 292294 209088 292350
rect 208768 292226 209088 292294
rect 208768 292170 208838 292226
rect 208894 292170 208962 292226
rect 209018 292170 209088 292226
rect 208768 292102 209088 292170
rect 208768 292046 208838 292102
rect 208894 292046 208962 292102
rect 209018 292046 209088 292102
rect 208768 291978 209088 292046
rect 208768 291922 208838 291978
rect 208894 291922 208962 291978
rect 209018 291922 209088 291978
rect 208768 291888 209088 291922
rect 239488 292350 239808 292384
rect 239488 292294 239558 292350
rect 239614 292294 239682 292350
rect 239738 292294 239808 292350
rect 239488 292226 239808 292294
rect 239488 292170 239558 292226
rect 239614 292170 239682 292226
rect 239738 292170 239808 292226
rect 239488 292102 239808 292170
rect 239488 292046 239558 292102
rect 239614 292046 239682 292102
rect 239738 292046 239808 292102
rect 239488 291978 239808 292046
rect 239488 291922 239558 291978
rect 239614 291922 239682 291978
rect 239738 291922 239808 291978
rect 239488 291888 239808 291922
rect 270208 292350 270528 292384
rect 270208 292294 270278 292350
rect 270334 292294 270402 292350
rect 270458 292294 270528 292350
rect 270208 292226 270528 292294
rect 270208 292170 270278 292226
rect 270334 292170 270402 292226
rect 270458 292170 270528 292226
rect 270208 292102 270528 292170
rect 270208 292046 270278 292102
rect 270334 292046 270402 292102
rect 270458 292046 270528 292102
rect 270208 291978 270528 292046
rect 270208 291922 270278 291978
rect 270334 291922 270402 291978
rect 270458 291922 270528 291978
rect 270208 291888 270528 291922
rect 300928 292350 301248 292384
rect 300928 292294 300998 292350
rect 301054 292294 301122 292350
rect 301178 292294 301248 292350
rect 300928 292226 301248 292294
rect 300928 292170 300998 292226
rect 301054 292170 301122 292226
rect 301178 292170 301248 292226
rect 300928 292102 301248 292170
rect 300928 292046 300998 292102
rect 301054 292046 301122 292102
rect 301178 292046 301248 292102
rect 300928 291978 301248 292046
rect 300928 291922 300998 291978
rect 301054 291922 301122 291978
rect 301178 291922 301248 291978
rect 300928 291888 301248 291922
rect 331648 292350 331968 292384
rect 331648 292294 331718 292350
rect 331774 292294 331842 292350
rect 331898 292294 331968 292350
rect 331648 292226 331968 292294
rect 331648 292170 331718 292226
rect 331774 292170 331842 292226
rect 331898 292170 331968 292226
rect 331648 292102 331968 292170
rect 331648 292046 331718 292102
rect 331774 292046 331842 292102
rect 331898 292046 331968 292102
rect 331648 291978 331968 292046
rect 331648 291922 331718 291978
rect 331774 291922 331842 291978
rect 331898 291922 331968 291978
rect 331648 291888 331968 291922
rect 362368 292350 362688 292384
rect 362368 292294 362438 292350
rect 362494 292294 362562 292350
rect 362618 292294 362688 292350
rect 362368 292226 362688 292294
rect 362368 292170 362438 292226
rect 362494 292170 362562 292226
rect 362618 292170 362688 292226
rect 362368 292102 362688 292170
rect 362368 292046 362438 292102
rect 362494 292046 362562 292102
rect 362618 292046 362688 292102
rect 362368 291978 362688 292046
rect 362368 291922 362438 291978
rect 362494 291922 362562 291978
rect 362618 291922 362688 291978
rect 362368 291888 362688 291922
rect 393088 292350 393408 292384
rect 393088 292294 393158 292350
rect 393214 292294 393282 292350
rect 393338 292294 393408 292350
rect 393088 292226 393408 292294
rect 393088 292170 393158 292226
rect 393214 292170 393282 292226
rect 393338 292170 393408 292226
rect 393088 292102 393408 292170
rect 393088 292046 393158 292102
rect 393214 292046 393282 292102
rect 393338 292046 393408 292102
rect 393088 291978 393408 292046
rect 393088 291922 393158 291978
rect 393214 291922 393282 291978
rect 393338 291922 393408 291978
rect 393088 291888 393408 291922
rect 423808 292350 424128 292384
rect 423808 292294 423878 292350
rect 423934 292294 424002 292350
rect 424058 292294 424128 292350
rect 423808 292226 424128 292294
rect 423808 292170 423878 292226
rect 423934 292170 424002 292226
rect 424058 292170 424128 292226
rect 423808 292102 424128 292170
rect 423808 292046 423878 292102
rect 423934 292046 424002 292102
rect 424058 292046 424128 292102
rect 423808 291978 424128 292046
rect 423808 291922 423878 291978
rect 423934 291922 424002 291978
rect 424058 291922 424128 291978
rect 423808 291888 424128 291922
rect 454528 292350 454848 292384
rect 454528 292294 454598 292350
rect 454654 292294 454722 292350
rect 454778 292294 454848 292350
rect 454528 292226 454848 292294
rect 454528 292170 454598 292226
rect 454654 292170 454722 292226
rect 454778 292170 454848 292226
rect 454528 292102 454848 292170
rect 454528 292046 454598 292102
rect 454654 292046 454722 292102
rect 454778 292046 454848 292102
rect 454528 291978 454848 292046
rect 454528 291922 454598 291978
rect 454654 291922 454722 291978
rect 454778 291922 454848 291978
rect 454528 291888 454848 291922
rect 485248 292350 485568 292384
rect 485248 292294 485318 292350
rect 485374 292294 485442 292350
rect 485498 292294 485568 292350
rect 485248 292226 485568 292294
rect 485248 292170 485318 292226
rect 485374 292170 485442 292226
rect 485498 292170 485568 292226
rect 485248 292102 485568 292170
rect 485248 292046 485318 292102
rect 485374 292046 485442 292102
rect 485498 292046 485568 292102
rect 485248 291978 485568 292046
rect 485248 291922 485318 291978
rect 485374 291922 485442 291978
rect 485498 291922 485568 291978
rect 485248 291888 485568 291922
rect 515968 292350 516288 292384
rect 515968 292294 516038 292350
rect 516094 292294 516162 292350
rect 516218 292294 516288 292350
rect 515968 292226 516288 292294
rect 515968 292170 516038 292226
rect 516094 292170 516162 292226
rect 516218 292170 516288 292226
rect 515968 292102 516288 292170
rect 515968 292046 516038 292102
rect 516094 292046 516162 292102
rect 516218 292046 516288 292102
rect 515968 291978 516288 292046
rect 515968 291922 516038 291978
rect 516094 291922 516162 291978
rect 516218 291922 516288 291978
rect 515968 291888 516288 291922
rect 525154 292350 525774 309922
rect 525154 292294 525250 292350
rect 525306 292294 525374 292350
rect 525430 292294 525498 292350
rect 525554 292294 525622 292350
rect 525678 292294 525774 292350
rect 525154 292226 525774 292294
rect 525154 292170 525250 292226
rect 525306 292170 525374 292226
rect 525430 292170 525498 292226
rect 525554 292170 525622 292226
rect 525678 292170 525774 292226
rect 525154 292102 525774 292170
rect 525154 292046 525250 292102
rect 525306 292046 525374 292102
rect 525430 292046 525498 292102
rect 525554 292046 525622 292102
rect 525678 292046 525774 292102
rect 525154 291978 525774 292046
rect 525154 291922 525250 291978
rect 525306 291922 525374 291978
rect 525430 291922 525498 291978
rect 525554 291922 525622 291978
rect 525678 291922 525774 291978
rect 6874 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 7494 280350
rect 6874 280226 7494 280294
rect 6874 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 7494 280226
rect 6874 280102 7494 280170
rect 6874 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 7494 280102
rect 6874 279978 7494 280046
rect 6874 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 7494 279978
rect 6874 262350 7494 279922
rect 39808 280350 40128 280384
rect 39808 280294 39878 280350
rect 39934 280294 40002 280350
rect 40058 280294 40128 280350
rect 39808 280226 40128 280294
rect 39808 280170 39878 280226
rect 39934 280170 40002 280226
rect 40058 280170 40128 280226
rect 39808 280102 40128 280170
rect 39808 280046 39878 280102
rect 39934 280046 40002 280102
rect 40058 280046 40128 280102
rect 39808 279978 40128 280046
rect 39808 279922 39878 279978
rect 39934 279922 40002 279978
rect 40058 279922 40128 279978
rect 39808 279888 40128 279922
rect 70528 280350 70848 280384
rect 70528 280294 70598 280350
rect 70654 280294 70722 280350
rect 70778 280294 70848 280350
rect 70528 280226 70848 280294
rect 70528 280170 70598 280226
rect 70654 280170 70722 280226
rect 70778 280170 70848 280226
rect 70528 280102 70848 280170
rect 70528 280046 70598 280102
rect 70654 280046 70722 280102
rect 70778 280046 70848 280102
rect 70528 279978 70848 280046
rect 70528 279922 70598 279978
rect 70654 279922 70722 279978
rect 70778 279922 70848 279978
rect 70528 279888 70848 279922
rect 101248 280350 101568 280384
rect 101248 280294 101318 280350
rect 101374 280294 101442 280350
rect 101498 280294 101568 280350
rect 101248 280226 101568 280294
rect 101248 280170 101318 280226
rect 101374 280170 101442 280226
rect 101498 280170 101568 280226
rect 101248 280102 101568 280170
rect 101248 280046 101318 280102
rect 101374 280046 101442 280102
rect 101498 280046 101568 280102
rect 101248 279978 101568 280046
rect 101248 279922 101318 279978
rect 101374 279922 101442 279978
rect 101498 279922 101568 279978
rect 101248 279888 101568 279922
rect 131968 280350 132288 280384
rect 131968 280294 132038 280350
rect 132094 280294 132162 280350
rect 132218 280294 132288 280350
rect 131968 280226 132288 280294
rect 131968 280170 132038 280226
rect 132094 280170 132162 280226
rect 132218 280170 132288 280226
rect 131968 280102 132288 280170
rect 131968 280046 132038 280102
rect 132094 280046 132162 280102
rect 132218 280046 132288 280102
rect 131968 279978 132288 280046
rect 131968 279922 132038 279978
rect 132094 279922 132162 279978
rect 132218 279922 132288 279978
rect 131968 279888 132288 279922
rect 162688 280350 163008 280384
rect 162688 280294 162758 280350
rect 162814 280294 162882 280350
rect 162938 280294 163008 280350
rect 162688 280226 163008 280294
rect 162688 280170 162758 280226
rect 162814 280170 162882 280226
rect 162938 280170 163008 280226
rect 162688 280102 163008 280170
rect 162688 280046 162758 280102
rect 162814 280046 162882 280102
rect 162938 280046 163008 280102
rect 162688 279978 163008 280046
rect 162688 279922 162758 279978
rect 162814 279922 162882 279978
rect 162938 279922 163008 279978
rect 162688 279888 163008 279922
rect 193408 280350 193728 280384
rect 193408 280294 193478 280350
rect 193534 280294 193602 280350
rect 193658 280294 193728 280350
rect 193408 280226 193728 280294
rect 193408 280170 193478 280226
rect 193534 280170 193602 280226
rect 193658 280170 193728 280226
rect 193408 280102 193728 280170
rect 193408 280046 193478 280102
rect 193534 280046 193602 280102
rect 193658 280046 193728 280102
rect 193408 279978 193728 280046
rect 193408 279922 193478 279978
rect 193534 279922 193602 279978
rect 193658 279922 193728 279978
rect 193408 279888 193728 279922
rect 224128 280350 224448 280384
rect 224128 280294 224198 280350
rect 224254 280294 224322 280350
rect 224378 280294 224448 280350
rect 224128 280226 224448 280294
rect 224128 280170 224198 280226
rect 224254 280170 224322 280226
rect 224378 280170 224448 280226
rect 224128 280102 224448 280170
rect 224128 280046 224198 280102
rect 224254 280046 224322 280102
rect 224378 280046 224448 280102
rect 224128 279978 224448 280046
rect 224128 279922 224198 279978
rect 224254 279922 224322 279978
rect 224378 279922 224448 279978
rect 224128 279888 224448 279922
rect 254848 280350 255168 280384
rect 254848 280294 254918 280350
rect 254974 280294 255042 280350
rect 255098 280294 255168 280350
rect 254848 280226 255168 280294
rect 254848 280170 254918 280226
rect 254974 280170 255042 280226
rect 255098 280170 255168 280226
rect 254848 280102 255168 280170
rect 254848 280046 254918 280102
rect 254974 280046 255042 280102
rect 255098 280046 255168 280102
rect 254848 279978 255168 280046
rect 254848 279922 254918 279978
rect 254974 279922 255042 279978
rect 255098 279922 255168 279978
rect 254848 279888 255168 279922
rect 285568 280350 285888 280384
rect 285568 280294 285638 280350
rect 285694 280294 285762 280350
rect 285818 280294 285888 280350
rect 285568 280226 285888 280294
rect 285568 280170 285638 280226
rect 285694 280170 285762 280226
rect 285818 280170 285888 280226
rect 285568 280102 285888 280170
rect 285568 280046 285638 280102
rect 285694 280046 285762 280102
rect 285818 280046 285888 280102
rect 285568 279978 285888 280046
rect 285568 279922 285638 279978
rect 285694 279922 285762 279978
rect 285818 279922 285888 279978
rect 285568 279888 285888 279922
rect 316288 280350 316608 280384
rect 316288 280294 316358 280350
rect 316414 280294 316482 280350
rect 316538 280294 316608 280350
rect 316288 280226 316608 280294
rect 316288 280170 316358 280226
rect 316414 280170 316482 280226
rect 316538 280170 316608 280226
rect 316288 280102 316608 280170
rect 316288 280046 316358 280102
rect 316414 280046 316482 280102
rect 316538 280046 316608 280102
rect 316288 279978 316608 280046
rect 316288 279922 316358 279978
rect 316414 279922 316482 279978
rect 316538 279922 316608 279978
rect 316288 279888 316608 279922
rect 347008 280350 347328 280384
rect 347008 280294 347078 280350
rect 347134 280294 347202 280350
rect 347258 280294 347328 280350
rect 347008 280226 347328 280294
rect 347008 280170 347078 280226
rect 347134 280170 347202 280226
rect 347258 280170 347328 280226
rect 347008 280102 347328 280170
rect 347008 280046 347078 280102
rect 347134 280046 347202 280102
rect 347258 280046 347328 280102
rect 347008 279978 347328 280046
rect 347008 279922 347078 279978
rect 347134 279922 347202 279978
rect 347258 279922 347328 279978
rect 347008 279888 347328 279922
rect 377728 280350 378048 280384
rect 377728 280294 377798 280350
rect 377854 280294 377922 280350
rect 377978 280294 378048 280350
rect 377728 280226 378048 280294
rect 377728 280170 377798 280226
rect 377854 280170 377922 280226
rect 377978 280170 378048 280226
rect 377728 280102 378048 280170
rect 377728 280046 377798 280102
rect 377854 280046 377922 280102
rect 377978 280046 378048 280102
rect 377728 279978 378048 280046
rect 377728 279922 377798 279978
rect 377854 279922 377922 279978
rect 377978 279922 378048 279978
rect 377728 279888 378048 279922
rect 408448 280350 408768 280384
rect 408448 280294 408518 280350
rect 408574 280294 408642 280350
rect 408698 280294 408768 280350
rect 408448 280226 408768 280294
rect 408448 280170 408518 280226
rect 408574 280170 408642 280226
rect 408698 280170 408768 280226
rect 408448 280102 408768 280170
rect 408448 280046 408518 280102
rect 408574 280046 408642 280102
rect 408698 280046 408768 280102
rect 408448 279978 408768 280046
rect 408448 279922 408518 279978
rect 408574 279922 408642 279978
rect 408698 279922 408768 279978
rect 408448 279888 408768 279922
rect 439168 280350 439488 280384
rect 439168 280294 439238 280350
rect 439294 280294 439362 280350
rect 439418 280294 439488 280350
rect 439168 280226 439488 280294
rect 439168 280170 439238 280226
rect 439294 280170 439362 280226
rect 439418 280170 439488 280226
rect 439168 280102 439488 280170
rect 439168 280046 439238 280102
rect 439294 280046 439362 280102
rect 439418 280046 439488 280102
rect 439168 279978 439488 280046
rect 439168 279922 439238 279978
rect 439294 279922 439362 279978
rect 439418 279922 439488 279978
rect 439168 279888 439488 279922
rect 469888 280350 470208 280384
rect 469888 280294 469958 280350
rect 470014 280294 470082 280350
rect 470138 280294 470208 280350
rect 469888 280226 470208 280294
rect 469888 280170 469958 280226
rect 470014 280170 470082 280226
rect 470138 280170 470208 280226
rect 469888 280102 470208 280170
rect 469888 280046 469958 280102
rect 470014 280046 470082 280102
rect 470138 280046 470208 280102
rect 469888 279978 470208 280046
rect 469888 279922 469958 279978
rect 470014 279922 470082 279978
rect 470138 279922 470208 279978
rect 469888 279888 470208 279922
rect 500608 280350 500928 280384
rect 500608 280294 500678 280350
rect 500734 280294 500802 280350
rect 500858 280294 500928 280350
rect 500608 280226 500928 280294
rect 500608 280170 500678 280226
rect 500734 280170 500802 280226
rect 500858 280170 500928 280226
rect 500608 280102 500928 280170
rect 500608 280046 500678 280102
rect 500734 280046 500802 280102
rect 500858 280046 500928 280102
rect 500608 279978 500928 280046
rect 500608 279922 500678 279978
rect 500734 279922 500802 279978
rect 500858 279922 500928 279978
rect 500608 279888 500928 279922
rect 24448 274350 24768 274384
rect 24448 274294 24518 274350
rect 24574 274294 24642 274350
rect 24698 274294 24768 274350
rect 24448 274226 24768 274294
rect 24448 274170 24518 274226
rect 24574 274170 24642 274226
rect 24698 274170 24768 274226
rect 24448 274102 24768 274170
rect 24448 274046 24518 274102
rect 24574 274046 24642 274102
rect 24698 274046 24768 274102
rect 24448 273978 24768 274046
rect 24448 273922 24518 273978
rect 24574 273922 24642 273978
rect 24698 273922 24768 273978
rect 24448 273888 24768 273922
rect 55168 274350 55488 274384
rect 55168 274294 55238 274350
rect 55294 274294 55362 274350
rect 55418 274294 55488 274350
rect 55168 274226 55488 274294
rect 55168 274170 55238 274226
rect 55294 274170 55362 274226
rect 55418 274170 55488 274226
rect 55168 274102 55488 274170
rect 55168 274046 55238 274102
rect 55294 274046 55362 274102
rect 55418 274046 55488 274102
rect 55168 273978 55488 274046
rect 55168 273922 55238 273978
rect 55294 273922 55362 273978
rect 55418 273922 55488 273978
rect 55168 273888 55488 273922
rect 85888 274350 86208 274384
rect 85888 274294 85958 274350
rect 86014 274294 86082 274350
rect 86138 274294 86208 274350
rect 85888 274226 86208 274294
rect 85888 274170 85958 274226
rect 86014 274170 86082 274226
rect 86138 274170 86208 274226
rect 85888 274102 86208 274170
rect 85888 274046 85958 274102
rect 86014 274046 86082 274102
rect 86138 274046 86208 274102
rect 85888 273978 86208 274046
rect 85888 273922 85958 273978
rect 86014 273922 86082 273978
rect 86138 273922 86208 273978
rect 85888 273888 86208 273922
rect 116608 274350 116928 274384
rect 116608 274294 116678 274350
rect 116734 274294 116802 274350
rect 116858 274294 116928 274350
rect 116608 274226 116928 274294
rect 116608 274170 116678 274226
rect 116734 274170 116802 274226
rect 116858 274170 116928 274226
rect 116608 274102 116928 274170
rect 116608 274046 116678 274102
rect 116734 274046 116802 274102
rect 116858 274046 116928 274102
rect 116608 273978 116928 274046
rect 116608 273922 116678 273978
rect 116734 273922 116802 273978
rect 116858 273922 116928 273978
rect 116608 273888 116928 273922
rect 147328 274350 147648 274384
rect 147328 274294 147398 274350
rect 147454 274294 147522 274350
rect 147578 274294 147648 274350
rect 147328 274226 147648 274294
rect 147328 274170 147398 274226
rect 147454 274170 147522 274226
rect 147578 274170 147648 274226
rect 147328 274102 147648 274170
rect 147328 274046 147398 274102
rect 147454 274046 147522 274102
rect 147578 274046 147648 274102
rect 147328 273978 147648 274046
rect 147328 273922 147398 273978
rect 147454 273922 147522 273978
rect 147578 273922 147648 273978
rect 147328 273888 147648 273922
rect 178048 274350 178368 274384
rect 178048 274294 178118 274350
rect 178174 274294 178242 274350
rect 178298 274294 178368 274350
rect 178048 274226 178368 274294
rect 178048 274170 178118 274226
rect 178174 274170 178242 274226
rect 178298 274170 178368 274226
rect 178048 274102 178368 274170
rect 178048 274046 178118 274102
rect 178174 274046 178242 274102
rect 178298 274046 178368 274102
rect 178048 273978 178368 274046
rect 178048 273922 178118 273978
rect 178174 273922 178242 273978
rect 178298 273922 178368 273978
rect 178048 273888 178368 273922
rect 208768 274350 209088 274384
rect 208768 274294 208838 274350
rect 208894 274294 208962 274350
rect 209018 274294 209088 274350
rect 208768 274226 209088 274294
rect 208768 274170 208838 274226
rect 208894 274170 208962 274226
rect 209018 274170 209088 274226
rect 208768 274102 209088 274170
rect 208768 274046 208838 274102
rect 208894 274046 208962 274102
rect 209018 274046 209088 274102
rect 208768 273978 209088 274046
rect 208768 273922 208838 273978
rect 208894 273922 208962 273978
rect 209018 273922 209088 273978
rect 208768 273888 209088 273922
rect 239488 274350 239808 274384
rect 239488 274294 239558 274350
rect 239614 274294 239682 274350
rect 239738 274294 239808 274350
rect 239488 274226 239808 274294
rect 239488 274170 239558 274226
rect 239614 274170 239682 274226
rect 239738 274170 239808 274226
rect 239488 274102 239808 274170
rect 239488 274046 239558 274102
rect 239614 274046 239682 274102
rect 239738 274046 239808 274102
rect 239488 273978 239808 274046
rect 239488 273922 239558 273978
rect 239614 273922 239682 273978
rect 239738 273922 239808 273978
rect 239488 273888 239808 273922
rect 270208 274350 270528 274384
rect 270208 274294 270278 274350
rect 270334 274294 270402 274350
rect 270458 274294 270528 274350
rect 270208 274226 270528 274294
rect 270208 274170 270278 274226
rect 270334 274170 270402 274226
rect 270458 274170 270528 274226
rect 270208 274102 270528 274170
rect 270208 274046 270278 274102
rect 270334 274046 270402 274102
rect 270458 274046 270528 274102
rect 270208 273978 270528 274046
rect 270208 273922 270278 273978
rect 270334 273922 270402 273978
rect 270458 273922 270528 273978
rect 270208 273888 270528 273922
rect 300928 274350 301248 274384
rect 300928 274294 300998 274350
rect 301054 274294 301122 274350
rect 301178 274294 301248 274350
rect 300928 274226 301248 274294
rect 300928 274170 300998 274226
rect 301054 274170 301122 274226
rect 301178 274170 301248 274226
rect 300928 274102 301248 274170
rect 300928 274046 300998 274102
rect 301054 274046 301122 274102
rect 301178 274046 301248 274102
rect 300928 273978 301248 274046
rect 300928 273922 300998 273978
rect 301054 273922 301122 273978
rect 301178 273922 301248 273978
rect 300928 273888 301248 273922
rect 331648 274350 331968 274384
rect 331648 274294 331718 274350
rect 331774 274294 331842 274350
rect 331898 274294 331968 274350
rect 331648 274226 331968 274294
rect 331648 274170 331718 274226
rect 331774 274170 331842 274226
rect 331898 274170 331968 274226
rect 331648 274102 331968 274170
rect 331648 274046 331718 274102
rect 331774 274046 331842 274102
rect 331898 274046 331968 274102
rect 331648 273978 331968 274046
rect 331648 273922 331718 273978
rect 331774 273922 331842 273978
rect 331898 273922 331968 273978
rect 331648 273888 331968 273922
rect 362368 274350 362688 274384
rect 362368 274294 362438 274350
rect 362494 274294 362562 274350
rect 362618 274294 362688 274350
rect 362368 274226 362688 274294
rect 362368 274170 362438 274226
rect 362494 274170 362562 274226
rect 362618 274170 362688 274226
rect 362368 274102 362688 274170
rect 362368 274046 362438 274102
rect 362494 274046 362562 274102
rect 362618 274046 362688 274102
rect 362368 273978 362688 274046
rect 362368 273922 362438 273978
rect 362494 273922 362562 273978
rect 362618 273922 362688 273978
rect 362368 273888 362688 273922
rect 393088 274350 393408 274384
rect 393088 274294 393158 274350
rect 393214 274294 393282 274350
rect 393338 274294 393408 274350
rect 393088 274226 393408 274294
rect 393088 274170 393158 274226
rect 393214 274170 393282 274226
rect 393338 274170 393408 274226
rect 393088 274102 393408 274170
rect 393088 274046 393158 274102
rect 393214 274046 393282 274102
rect 393338 274046 393408 274102
rect 393088 273978 393408 274046
rect 393088 273922 393158 273978
rect 393214 273922 393282 273978
rect 393338 273922 393408 273978
rect 393088 273888 393408 273922
rect 423808 274350 424128 274384
rect 423808 274294 423878 274350
rect 423934 274294 424002 274350
rect 424058 274294 424128 274350
rect 423808 274226 424128 274294
rect 423808 274170 423878 274226
rect 423934 274170 424002 274226
rect 424058 274170 424128 274226
rect 423808 274102 424128 274170
rect 423808 274046 423878 274102
rect 423934 274046 424002 274102
rect 424058 274046 424128 274102
rect 423808 273978 424128 274046
rect 423808 273922 423878 273978
rect 423934 273922 424002 273978
rect 424058 273922 424128 273978
rect 423808 273888 424128 273922
rect 454528 274350 454848 274384
rect 454528 274294 454598 274350
rect 454654 274294 454722 274350
rect 454778 274294 454848 274350
rect 454528 274226 454848 274294
rect 454528 274170 454598 274226
rect 454654 274170 454722 274226
rect 454778 274170 454848 274226
rect 454528 274102 454848 274170
rect 454528 274046 454598 274102
rect 454654 274046 454722 274102
rect 454778 274046 454848 274102
rect 454528 273978 454848 274046
rect 454528 273922 454598 273978
rect 454654 273922 454722 273978
rect 454778 273922 454848 273978
rect 454528 273888 454848 273922
rect 485248 274350 485568 274384
rect 485248 274294 485318 274350
rect 485374 274294 485442 274350
rect 485498 274294 485568 274350
rect 485248 274226 485568 274294
rect 485248 274170 485318 274226
rect 485374 274170 485442 274226
rect 485498 274170 485568 274226
rect 485248 274102 485568 274170
rect 485248 274046 485318 274102
rect 485374 274046 485442 274102
rect 485498 274046 485568 274102
rect 485248 273978 485568 274046
rect 485248 273922 485318 273978
rect 485374 273922 485442 273978
rect 485498 273922 485568 273978
rect 485248 273888 485568 273922
rect 515968 274350 516288 274384
rect 515968 274294 516038 274350
rect 516094 274294 516162 274350
rect 516218 274294 516288 274350
rect 515968 274226 516288 274294
rect 515968 274170 516038 274226
rect 516094 274170 516162 274226
rect 516218 274170 516288 274226
rect 515968 274102 516288 274170
rect 515968 274046 516038 274102
rect 516094 274046 516162 274102
rect 516218 274046 516288 274102
rect 515968 273978 516288 274046
rect 515968 273922 516038 273978
rect 516094 273922 516162 273978
rect 516218 273922 516288 273978
rect 515968 273888 516288 273922
rect 525154 274350 525774 291922
rect 525154 274294 525250 274350
rect 525306 274294 525374 274350
rect 525430 274294 525498 274350
rect 525554 274294 525622 274350
rect 525678 274294 525774 274350
rect 525154 274226 525774 274294
rect 525154 274170 525250 274226
rect 525306 274170 525374 274226
rect 525430 274170 525498 274226
rect 525554 274170 525622 274226
rect 525678 274170 525774 274226
rect 525154 274102 525774 274170
rect 525154 274046 525250 274102
rect 525306 274046 525374 274102
rect 525430 274046 525498 274102
rect 525554 274046 525622 274102
rect 525678 274046 525774 274102
rect 525154 273978 525774 274046
rect 525154 273922 525250 273978
rect 525306 273922 525374 273978
rect 525430 273922 525498 273978
rect 525554 273922 525622 273978
rect 525678 273922 525774 273978
rect 6874 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 7494 262350
rect 6874 262226 7494 262294
rect 6874 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 7494 262226
rect 6874 262102 7494 262170
rect 6874 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 7494 262102
rect 6874 261978 7494 262046
rect 6874 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 7494 261978
rect 6874 244350 7494 261922
rect 39808 262350 40128 262384
rect 39808 262294 39878 262350
rect 39934 262294 40002 262350
rect 40058 262294 40128 262350
rect 39808 262226 40128 262294
rect 39808 262170 39878 262226
rect 39934 262170 40002 262226
rect 40058 262170 40128 262226
rect 39808 262102 40128 262170
rect 39808 262046 39878 262102
rect 39934 262046 40002 262102
rect 40058 262046 40128 262102
rect 39808 261978 40128 262046
rect 39808 261922 39878 261978
rect 39934 261922 40002 261978
rect 40058 261922 40128 261978
rect 39808 261888 40128 261922
rect 70528 262350 70848 262384
rect 70528 262294 70598 262350
rect 70654 262294 70722 262350
rect 70778 262294 70848 262350
rect 70528 262226 70848 262294
rect 70528 262170 70598 262226
rect 70654 262170 70722 262226
rect 70778 262170 70848 262226
rect 70528 262102 70848 262170
rect 70528 262046 70598 262102
rect 70654 262046 70722 262102
rect 70778 262046 70848 262102
rect 70528 261978 70848 262046
rect 70528 261922 70598 261978
rect 70654 261922 70722 261978
rect 70778 261922 70848 261978
rect 70528 261888 70848 261922
rect 101248 262350 101568 262384
rect 101248 262294 101318 262350
rect 101374 262294 101442 262350
rect 101498 262294 101568 262350
rect 101248 262226 101568 262294
rect 101248 262170 101318 262226
rect 101374 262170 101442 262226
rect 101498 262170 101568 262226
rect 101248 262102 101568 262170
rect 101248 262046 101318 262102
rect 101374 262046 101442 262102
rect 101498 262046 101568 262102
rect 101248 261978 101568 262046
rect 101248 261922 101318 261978
rect 101374 261922 101442 261978
rect 101498 261922 101568 261978
rect 101248 261888 101568 261922
rect 131968 262350 132288 262384
rect 131968 262294 132038 262350
rect 132094 262294 132162 262350
rect 132218 262294 132288 262350
rect 131968 262226 132288 262294
rect 131968 262170 132038 262226
rect 132094 262170 132162 262226
rect 132218 262170 132288 262226
rect 131968 262102 132288 262170
rect 131968 262046 132038 262102
rect 132094 262046 132162 262102
rect 132218 262046 132288 262102
rect 131968 261978 132288 262046
rect 131968 261922 132038 261978
rect 132094 261922 132162 261978
rect 132218 261922 132288 261978
rect 131968 261888 132288 261922
rect 162688 262350 163008 262384
rect 162688 262294 162758 262350
rect 162814 262294 162882 262350
rect 162938 262294 163008 262350
rect 162688 262226 163008 262294
rect 162688 262170 162758 262226
rect 162814 262170 162882 262226
rect 162938 262170 163008 262226
rect 162688 262102 163008 262170
rect 162688 262046 162758 262102
rect 162814 262046 162882 262102
rect 162938 262046 163008 262102
rect 162688 261978 163008 262046
rect 162688 261922 162758 261978
rect 162814 261922 162882 261978
rect 162938 261922 163008 261978
rect 162688 261888 163008 261922
rect 193408 262350 193728 262384
rect 193408 262294 193478 262350
rect 193534 262294 193602 262350
rect 193658 262294 193728 262350
rect 193408 262226 193728 262294
rect 193408 262170 193478 262226
rect 193534 262170 193602 262226
rect 193658 262170 193728 262226
rect 193408 262102 193728 262170
rect 193408 262046 193478 262102
rect 193534 262046 193602 262102
rect 193658 262046 193728 262102
rect 193408 261978 193728 262046
rect 193408 261922 193478 261978
rect 193534 261922 193602 261978
rect 193658 261922 193728 261978
rect 193408 261888 193728 261922
rect 224128 262350 224448 262384
rect 224128 262294 224198 262350
rect 224254 262294 224322 262350
rect 224378 262294 224448 262350
rect 224128 262226 224448 262294
rect 224128 262170 224198 262226
rect 224254 262170 224322 262226
rect 224378 262170 224448 262226
rect 224128 262102 224448 262170
rect 224128 262046 224198 262102
rect 224254 262046 224322 262102
rect 224378 262046 224448 262102
rect 224128 261978 224448 262046
rect 224128 261922 224198 261978
rect 224254 261922 224322 261978
rect 224378 261922 224448 261978
rect 224128 261888 224448 261922
rect 254848 262350 255168 262384
rect 254848 262294 254918 262350
rect 254974 262294 255042 262350
rect 255098 262294 255168 262350
rect 254848 262226 255168 262294
rect 254848 262170 254918 262226
rect 254974 262170 255042 262226
rect 255098 262170 255168 262226
rect 254848 262102 255168 262170
rect 254848 262046 254918 262102
rect 254974 262046 255042 262102
rect 255098 262046 255168 262102
rect 254848 261978 255168 262046
rect 254848 261922 254918 261978
rect 254974 261922 255042 261978
rect 255098 261922 255168 261978
rect 254848 261888 255168 261922
rect 285568 262350 285888 262384
rect 285568 262294 285638 262350
rect 285694 262294 285762 262350
rect 285818 262294 285888 262350
rect 285568 262226 285888 262294
rect 285568 262170 285638 262226
rect 285694 262170 285762 262226
rect 285818 262170 285888 262226
rect 285568 262102 285888 262170
rect 285568 262046 285638 262102
rect 285694 262046 285762 262102
rect 285818 262046 285888 262102
rect 285568 261978 285888 262046
rect 285568 261922 285638 261978
rect 285694 261922 285762 261978
rect 285818 261922 285888 261978
rect 285568 261888 285888 261922
rect 316288 262350 316608 262384
rect 316288 262294 316358 262350
rect 316414 262294 316482 262350
rect 316538 262294 316608 262350
rect 316288 262226 316608 262294
rect 316288 262170 316358 262226
rect 316414 262170 316482 262226
rect 316538 262170 316608 262226
rect 316288 262102 316608 262170
rect 316288 262046 316358 262102
rect 316414 262046 316482 262102
rect 316538 262046 316608 262102
rect 316288 261978 316608 262046
rect 316288 261922 316358 261978
rect 316414 261922 316482 261978
rect 316538 261922 316608 261978
rect 316288 261888 316608 261922
rect 347008 262350 347328 262384
rect 347008 262294 347078 262350
rect 347134 262294 347202 262350
rect 347258 262294 347328 262350
rect 347008 262226 347328 262294
rect 347008 262170 347078 262226
rect 347134 262170 347202 262226
rect 347258 262170 347328 262226
rect 347008 262102 347328 262170
rect 347008 262046 347078 262102
rect 347134 262046 347202 262102
rect 347258 262046 347328 262102
rect 347008 261978 347328 262046
rect 347008 261922 347078 261978
rect 347134 261922 347202 261978
rect 347258 261922 347328 261978
rect 347008 261888 347328 261922
rect 377728 262350 378048 262384
rect 377728 262294 377798 262350
rect 377854 262294 377922 262350
rect 377978 262294 378048 262350
rect 377728 262226 378048 262294
rect 377728 262170 377798 262226
rect 377854 262170 377922 262226
rect 377978 262170 378048 262226
rect 377728 262102 378048 262170
rect 377728 262046 377798 262102
rect 377854 262046 377922 262102
rect 377978 262046 378048 262102
rect 377728 261978 378048 262046
rect 377728 261922 377798 261978
rect 377854 261922 377922 261978
rect 377978 261922 378048 261978
rect 377728 261888 378048 261922
rect 408448 262350 408768 262384
rect 408448 262294 408518 262350
rect 408574 262294 408642 262350
rect 408698 262294 408768 262350
rect 408448 262226 408768 262294
rect 408448 262170 408518 262226
rect 408574 262170 408642 262226
rect 408698 262170 408768 262226
rect 408448 262102 408768 262170
rect 408448 262046 408518 262102
rect 408574 262046 408642 262102
rect 408698 262046 408768 262102
rect 408448 261978 408768 262046
rect 408448 261922 408518 261978
rect 408574 261922 408642 261978
rect 408698 261922 408768 261978
rect 408448 261888 408768 261922
rect 439168 262350 439488 262384
rect 439168 262294 439238 262350
rect 439294 262294 439362 262350
rect 439418 262294 439488 262350
rect 439168 262226 439488 262294
rect 439168 262170 439238 262226
rect 439294 262170 439362 262226
rect 439418 262170 439488 262226
rect 439168 262102 439488 262170
rect 439168 262046 439238 262102
rect 439294 262046 439362 262102
rect 439418 262046 439488 262102
rect 439168 261978 439488 262046
rect 439168 261922 439238 261978
rect 439294 261922 439362 261978
rect 439418 261922 439488 261978
rect 439168 261888 439488 261922
rect 469888 262350 470208 262384
rect 469888 262294 469958 262350
rect 470014 262294 470082 262350
rect 470138 262294 470208 262350
rect 469888 262226 470208 262294
rect 469888 262170 469958 262226
rect 470014 262170 470082 262226
rect 470138 262170 470208 262226
rect 469888 262102 470208 262170
rect 469888 262046 469958 262102
rect 470014 262046 470082 262102
rect 470138 262046 470208 262102
rect 469888 261978 470208 262046
rect 469888 261922 469958 261978
rect 470014 261922 470082 261978
rect 470138 261922 470208 261978
rect 469888 261888 470208 261922
rect 500608 262350 500928 262384
rect 500608 262294 500678 262350
rect 500734 262294 500802 262350
rect 500858 262294 500928 262350
rect 500608 262226 500928 262294
rect 500608 262170 500678 262226
rect 500734 262170 500802 262226
rect 500858 262170 500928 262226
rect 500608 262102 500928 262170
rect 500608 262046 500678 262102
rect 500734 262046 500802 262102
rect 500858 262046 500928 262102
rect 500608 261978 500928 262046
rect 500608 261922 500678 261978
rect 500734 261922 500802 261978
rect 500858 261922 500928 261978
rect 500608 261888 500928 261922
rect 24448 256350 24768 256384
rect 24448 256294 24518 256350
rect 24574 256294 24642 256350
rect 24698 256294 24768 256350
rect 24448 256226 24768 256294
rect 24448 256170 24518 256226
rect 24574 256170 24642 256226
rect 24698 256170 24768 256226
rect 24448 256102 24768 256170
rect 24448 256046 24518 256102
rect 24574 256046 24642 256102
rect 24698 256046 24768 256102
rect 24448 255978 24768 256046
rect 24448 255922 24518 255978
rect 24574 255922 24642 255978
rect 24698 255922 24768 255978
rect 24448 255888 24768 255922
rect 55168 256350 55488 256384
rect 55168 256294 55238 256350
rect 55294 256294 55362 256350
rect 55418 256294 55488 256350
rect 55168 256226 55488 256294
rect 55168 256170 55238 256226
rect 55294 256170 55362 256226
rect 55418 256170 55488 256226
rect 55168 256102 55488 256170
rect 55168 256046 55238 256102
rect 55294 256046 55362 256102
rect 55418 256046 55488 256102
rect 55168 255978 55488 256046
rect 55168 255922 55238 255978
rect 55294 255922 55362 255978
rect 55418 255922 55488 255978
rect 55168 255888 55488 255922
rect 85888 256350 86208 256384
rect 85888 256294 85958 256350
rect 86014 256294 86082 256350
rect 86138 256294 86208 256350
rect 85888 256226 86208 256294
rect 85888 256170 85958 256226
rect 86014 256170 86082 256226
rect 86138 256170 86208 256226
rect 85888 256102 86208 256170
rect 85888 256046 85958 256102
rect 86014 256046 86082 256102
rect 86138 256046 86208 256102
rect 85888 255978 86208 256046
rect 85888 255922 85958 255978
rect 86014 255922 86082 255978
rect 86138 255922 86208 255978
rect 85888 255888 86208 255922
rect 116608 256350 116928 256384
rect 116608 256294 116678 256350
rect 116734 256294 116802 256350
rect 116858 256294 116928 256350
rect 116608 256226 116928 256294
rect 116608 256170 116678 256226
rect 116734 256170 116802 256226
rect 116858 256170 116928 256226
rect 116608 256102 116928 256170
rect 116608 256046 116678 256102
rect 116734 256046 116802 256102
rect 116858 256046 116928 256102
rect 116608 255978 116928 256046
rect 116608 255922 116678 255978
rect 116734 255922 116802 255978
rect 116858 255922 116928 255978
rect 116608 255888 116928 255922
rect 147328 256350 147648 256384
rect 147328 256294 147398 256350
rect 147454 256294 147522 256350
rect 147578 256294 147648 256350
rect 147328 256226 147648 256294
rect 147328 256170 147398 256226
rect 147454 256170 147522 256226
rect 147578 256170 147648 256226
rect 147328 256102 147648 256170
rect 147328 256046 147398 256102
rect 147454 256046 147522 256102
rect 147578 256046 147648 256102
rect 147328 255978 147648 256046
rect 147328 255922 147398 255978
rect 147454 255922 147522 255978
rect 147578 255922 147648 255978
rect 147328 255888 147648 255922
rect 178048 256350 178368 256384
rect 178048 256294 178118 256350
rect 178174 256294 178242 256350
rect 178298 256294 178368 256350
rect 178048 256226 178368 256294
rect 178048 256170 178118 256226
rect 178174 256170 178242 256226
rect 178298 256170 178368 256226
rect 178048 256102 178368 256170
rect 178048 256046 178118 256102
rect 178174 256046 178242 256102
rect 178298 256046 178368 256102
rect 178048 255978 178368 256046
rect 178048 255922 178118 255978
rect 178174 255922 178242 255978
rect 178298 255922 178368 255978
rect 178048 255888 178368 255922
rect 208768 256350 209088 256384
rect 208768 256294 208838 256350
rect 208894 256294 208962 256350
rect 209018 256294 209088 256350
rect 208768 256226 209088 256294
rect 208768 256170 208838 256226
rect 208894 256170 208962 256226
rect 209018 256170 209088 256226
rect 208768 256102 209088 256170
rect 208768 256046 208838 256102
rect 208894 256046 208962 256102
rect 209018 256046 209088 256102
rect 208768 255978 209088 256046
rect 208768 255922 208838 255978
rect 208894 255922 208962 255978
rect 209018 255922 209088 255978
rect 208768 255888 209088 255922
rect 239488 256350 239808 256384
rect 239488 256294 239558 256350
rect 239614 256294 239682 256350
rect 239738 256294 239808 256350
rect 239488 256226 239808 256294
rect 239488 256170 239558 256226
rect 239614 256170 239682 256226
rect 239738 256170 239808 256226
rect 239488 256102 239808 256170
rect 239488 256046 239558 256102
rect 239614 256046 239682 256102
rect 239738 256046 239808 256102
rect 239488 255978 239808 256046
rect 239488 255922 239558 255978
rect 239614 255922 239682 255978
rect 239738 255922 239808 255978
rect 239488 255888 239808 255922
rect 270208 256350 270528 256384
rect 270208 256294 270278 256350
rect 270334 256294 270402 256350
rect 270458 256294 270528 256350
rect 270208 256226 270528 256294
rect 270208 256170 270278 256226
rect 270334 256170 270402 256226
rect 270458 256170 270528 256226
rect 270208 256102 270528 256170
rect 270208 256046 270278 256102
rect 270334 256046 270402 256102
rect 270458 256046 270528 256102
rect 270208 255978 270528 256046
rect 270208 255922 270278 255978
rect 270334 255922 270402 255978
rect 270458 255922 270528 255978
rect 270208 255888 270528 255922
rect 300928 256350 301248 256384
rect 300928 256294 300998 256350
rect 301054 256294 301122 256350
rect 301178 256294 301248 256350
rect 300928 256226 301248 256294
rect 300928 256170 300998 256226
rect 301054 256170 301122 256226
rect 301178 256170 301248 256226
rect 300928 256102 301248 256170
rect 300928 256046 300998 256102
rect 301054 256046 301122 256102
rect 301178 256046 301248 256102
rect 300928 255978 301248 256046
rect 300928 255922 300998 255978
rect 301054 255922 301122 255978
rect 301178 255922 301248 255978
rect 300928 255888 301248 255922
rect 331648 256350 331968 256384
rect 331648 256294 331718 256350
rect 331774 256294 331842 256350
rect 331898 256294 331968 256350
rect 331648 256226 331968 256294
rect 331648 256170 331718 256226
rect 331774 256170 331842 256226
rect 331898 256170 331968 256226
rect 331648 256102 331968 256170
rect 331648 256046 331718 256102
rect 331774 256046 331842 256102
rect 331898 256046 331968 256102
rect 331648 255978 331968 256046
rect 331648 255922 331718 255978
rect 331774 255922 331842 255978
rect 331898 255922 331968 255978
rect 331648 255888 331968 255922
rect 362368 256350 362688 256384
rect 362368 256294 362438 256350
rect 362494 256294 362562 256350
rect 362618 256294 362688 256350
rect 362368 256226 362688 256294
rect 362368 256170 362438 256226
rect 362494 256170 362562 256226
rect 362618 256170 362688 256226
rect 362368 256102 362688 256170
rect 362368 256046 362438 256102
rect 362494 256046 362562 256102
rect 362618 256046 362688 256102
rect 362368 255978 362688 256046
rect 362368 255922 362438 255978
rect 362494 255922 362562 255978
rect 362618 255922 362688 255978
rect 362368 255888 362688 255922
rect 393088 256350 393408 256384
rect 393088 256294 393158 256350
rect 393214 256294 393282 256350
rect 393338 256294 393408 256350
rect 393088 256226 393408 256294
rect 393088 256170 393158 256226
rect 393214 256170 393282 256226
rect 393338 256170 393408 256226
rect 393088 256102 393408 256170
rect 393088 256046 393158 256102
rect 393214 256046 393282 256102
rect 393338 256046 393408 256102
rect 393088 255978 393408 256046
rect 393088 255922 393158 255978
rect 393214 255922 393282 255978
rect 393338 255922 393408 255978
rect 393088 255888 393408 255922
rect 423808 256350 424128 256384
rect 423808 256294 423878 256350
rect 423934 256294 424002 256350
rect 424058 256294 424128 256350
rect 423808 256226 424128 256294
rect 423808 256170 423878 256226
rect 423934 256170 424002 256226
rect 424058 256170 424128 256226
rect 423808 256102 424128 256170
rect 423808 256046 423878 256102
rect 423934 256046 424002 256102
rect 424058 256046 424128 256102
rect 423808 255978 424128 256046
rect 423808 255922 423878 255978
rect 423934 255922 424002 255978
rect 424058 255922 424128 255978
rect 423808 255888 424128 255922
rect 454528 256350 454848 256384
rect 454528 256294 454598 256350
rect 454654 256294 454722 256350
rect 454778 256294 454848 256350
rect 454528 256226 454848 256294
rect 454528 256170 454598 256226
rect 454654 256170 454722 256226
rect 454778 256170 454848 256226
rect 454528 256102 454848 256170
rect 454528 256046 454598 256102
rect 454654 256046 454722 256102
rect 454778 256046 454848 256102
rect 454528 255978 454848 256046
rect 454528 255922 454598 255978
rect 454654 255922 454722 255978
rect 454778 255922 454848 255978
rect 454528 255888 454848 255922
rect 485248 256350 485568 256384
rect 485248 256294 485318 256350
rect 485374 256294 485442 256350
rect 485498 256294 485568 256350
rect 485248 256226 485568 256294
rect 485248 256170 485318 256226
rect 485374 256170 485442 256226
rect 485498 256170 485568 256226
rect 485248 256102 485568 256170
rect 485248 256046 485318 256102
rect 485374 256046 485442 256102
rect 485498 256046 485568 256102
rect 485248 255978 485568 256046
rect 485248 255922 485318 255978
rect 485374 255922 485442 255978
rect 485498 255922 485568 255978
rect 485248 255888 485568 255922
rect 515968 256350 516288 256384
rect 515968 256294 516038 256350
rect 516094 256294 516162 256350
rect 516218 256294 516288 256350
rect 515968 256226 516288 256294
rect 515968 256170 516038 256226
rect 516094 256170 516162 256226
rect 516218 256170 516288 256226
rect 515968 256102 516288 256170
rect 515968 256046 516038 256102
rect 516094 256046 516162 256102
rect 516218 256046 516288 256102
rect 515968 255978 516288 256046
rect 515968 255922 516038 255978
rect 516094 255922 516162 255978
rect 516218 255922 516288 255978
rect 515968 255888 516288 255922
rect 525154 256350 525774 273922
rect 525154 256294 525250 256350
rect 525306 256294 525374 256350
rect 525430 256294 525498 256350
rect 525554 256294 525622 256350
rect 525678 256294 525774 256350
rect 525154 256226 525774 256294
rect 525154 256170 525250 256226
rect 525306 256170 525374 256226
rect 525430 256170 525498 256226
rect 525554 256170 525622 256226
rect 525678 256170 525774 256226
rect 525154 256102 525774 256170
rect 525154 256046 525250 256102
rect 525306 256046 525374 256102
rect 525430 256046 525498 256102
rect 525554 256046 525622 256102
rect 525678 256046 525774 256102
rect 525154 255978 525774 256046
rect 525154 255922 525250 255978
rect 525306 255922 525374 255978
rect 525430 255922 525498 255978
rect 525554 255922 525622 255978
rect 525678 255922 525774 255978
rect 6874 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 7494 244350
rect 6874 244226 7494 244294
rect 6874 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 7494 244226
rect 6874 244102 7494 244170
rect 6874 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 7494 244102
rect 6874 243978 7494 244046
rect 6874 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 7494 243978
rect 6874 226350 7494 243922
rect 39808 244350 40128 244384
rect 39808 244294 39878 244350
rect 39934 244294 40002 244350
rect 40058 244294 40128 244350
rect 39808 244226 40128 244294
rect 39808 244170 39878 244226
rect 39934 244170 40002 244226
rect 40058 244170 40128 244226
rect 39808 244102 40128 244170
rect 39808 244046 39878 244102
rect 39934 244046 40002 244102
rect 40058 244046 40128 244102
rect 39808 243978 40128 244046
rect 39808 243922 39878 243978
rect 39934 243922 40002 243978
rect 40058 243922 40128 243978
rect 39808 243888 40128 243922
rect 70528 244350 70848 244384
rect 70528 244294 70598 244350
rect 70654 244294 70722 244350
rect 70778 244294 70848 244350
rect 70528 244226 70848 244294
rect 70528 244170 70598 244226
rect 70654 244170 70722 244226
rect 70778 244170 70848 244226
rect 70528 244102 70848 244170
rect 70528 244046 70598 244102
rect 70654 244046 70722 244102
rect 70778 244046 70848 244102
rect 70528 243978 70848 244046
rect 70528 243922 70598 243978
rect 70654 243922 70722 243978
rect 70778 243922 70848 243978
rect 70528 243888 70848 243922
rect 101248 244350 101568 244384
rect 101248 244294 101318 244350
rect 101374 244294 101442 244350
rect 101498 244294 101568 244350
rect 101248 244226 101568 244294
rect 101248 244170 101318 244226
rect 101374 244170 101442 244226
rect 101498 244170 101568 244226
rect 101248 244102 101568 244170
rect 101248 244046 101318 244102
rect 101374 244046 101442 244102
rect 101498 244046 101568 244102
rect 101248 243978 101568 244046
rect 101248 243922 101318 243978
rect 101374 243922 101442 243978
rect 101498 243922 101568 243978
rect 101248 243888 101568 243922
rect 131968 244350 132288 244384
rect 131968 244294 132038 244350
rect 132094 244294 132162 244350
rect 132218 244294 132288 244350
rect 131968 244226 132288 244294
rect 131968 244170 132038 244226
rect 132094 244170 132162 244226
rect 132218 244170 132288 244226
rect 131968 244102 132288 244170
rect 131968 244046 132038 244102
rect 132094 244046 132162 244102
rect 132218 244046 132288 244102
rect 131968 243978 132288 244046
rect 131968 243922 132038 243978
rect 132094 243922 132162 243978
rect 132218 243922 132288 243978
rect 131968 243888 132288 243922
rect 162688 244350 163008 244384
rect 162688 244294 162758 244350
rect 162814 244294 162882 244350
rect 162938 244294 163008 244350
rect 162688 244226 163008 244294
rect 162688 244170 162758 244226
rect 162814 244170 162882 244226
rect 162938 244170 163008 244226
rect 162688 244102 163008 244170
rect 162688 244046 162758 244102
rect 162814 244046 162882 244102
rect 162938 244046 163008 244102
rect 162688 243978 163008 244046
rect 162688 243922 162758 243978
rect 162814 243922 162882 243978
rect 162938 243922 163008 243978
rect 162688 243888 163008 243922
rect 193408 244350 193728 244384
rect 193408 244294 193478 244350
rect 193534 244294 193602 244350
rect 193658 244294 193728 244350
rect 193408 244226 193728 244294
rect 193408 244170 193478 244226
rect 193534 244170 193602 244226
rect 193658 244170 193728 244226
rect 193408 244102 193728 244170
rect 193408 244046 193478 244102
rect 193534 244046 193602 244102
rect 193658 244046 193728 244102
rect 193408 243978 193728 244046
rect 193408 243922 193478 243978
rect 193534 243922 193602 243978
rect 193658 243922 193728 243978
rect 193408 243888 193728 243922
rect 224128 244350 224448 244384
rect 224128 244294 224198 244350
rect 224254 244294 224322 244350
rect 224378 244294 224448 244350
rect 224128 244226 224448 244294
rect 224128 244170 224198 244226
rect 224254 244170 224322 244226
rect 224378 244170 224448 244226
rect 224128 244102 224448 244170
rect 224128 244046 224198 244102
rect 224254 244046 224322 244102
rect 224378 244046 224448 244102
rect 224128 243978 224448 244046
rect 224128 243922 224198 243978
rect 224254 243922 224322 243978
rect 224378 243922 224448 243978
rect 224128 243888 224448 243922
rect 254848 244350 255168 244384
rect 254848 244294 254918 244350
rect 254974 244294 255042 244350
rect 255098 244294 255168 244350
rect 254848 244226 255168 244294
rect 254848 244170 254918 244226
rect 254974 244170 255042 244226
rect 255098 244170 255168 244226
rect 254848 244102 255168 244170
rect 254848 244046 254918 244102
rect 254974 244046 255042 244102
rect 255098 244046 255168 244102
rect 254848 243978 255168 244046
rect 254848 243922 254918 243978
rect 254974 243922 255042 243978
rect 255098 243922 255168 243978
rect 254848 243888 255168 243922
rect 285568 244350 285888 244384
rect 285568 244294 285638 244350
rect 285694 244294 285762 244350
rect 285818 244294 285888 244350
rect 285568 244226 285888 244294
rect 285568 244170 285638 244226
rect 285694 244170 285762 244226
rect 285818 244170 285888 244226
rect 285568 244102 285888 244170
rect 285568 244046 285638 244102
rect 285694 244046 285762 244102
rect 285818 244046 285888 244102
rect 285568 243978 285888 244046
rect 285568 243922 285638 243978
rect 285694 243922 285762 243978
rect 285818 243922 285888 243978
rect 285568 243888 285888 243922
rect 316288 244350 316608 244384
rect 316288 244294 316358 244350
rect 316414 244294 316482 244350
rect 316538 244294 316608 244350
rect 316288 244226 316608 244294
rect 316288 244170 316358 244226
rect 316414 244170 316482 244226
rect 316538 244170 316608 244226
rect 316288 244102 316608 244170
rect 316288 244046 316358 244102
rect 316414 244046 316482 244102
rect 316538 244046 316608 244102
rect 316288 243978 316608 244046
rect 316288 243922 316358 243978
rect 316414 243922 316482 243978
rect 316538 243922 316608 243978
rect 316288 243888 316608 243922
rect 347008 244350 347328 244384
rect 347008 244294 347078 244350
rect 347134 244294 347202 244350
rect 347258 244294 347328 244350
rect 347008 244226 347328 244294
rect 347008 244170 347078 244226
rect 347134 244170 347202 244226
rect 347258 244170 347328 244226
rect 347008 244102 347328 244170
rect 347008 244046 347078 244102
rect 347134 244046 347202 244102
rect 347258 244046 347328 244102
rect 347008 243978 347328 244046
rect 347008 243922 347078 243978
rect 347134 243922 347202 243978
rect 347258 243922 347328 243978
rect 347008 243888 347328 243922
rect 377728 244350 378048 244384
rect 377728 244294 377798 244350
rect 377854 244294 377922 244350
rect 377978 244294 378048 244350
rect 377728 244226 378048 244294
rect 377728 244170 377798 244226
rect 377854 244170 377922 244226
rect 377978 244170 378048 244226
rect 377728 244102 378048 244170
rect 377728 244046 377798 244102
rect 377854 244046 377922 244102
rect 377978 244046 378048 244102
rect 377728 243978 378048 244046
rect 377728 243922 377798 243978
rect 377854 243922 377922 243978
rect 377978 243922 378048 243978
rect 377728 243888 378048 243922
rect 408448 244350 408768 244384
rect 408448 244294 408518 244350
rect 408574 244294 408642 244350
rect 408698 244294 408768 244350
rect 408448 244226 408768 244294
rect 408448 244170 408518 244226
rect 408574 244170 408642 244226
rect 408698 244170 408768 244226
rect 408448 244102 408768 244170
rect 408448 244046 408518 244102
rect 408574 244046 408642 244102
rect 408698 244046 408768 244102
rect 408448 243978 408768 244046
rect 408448 243922 408518 243978
rect 408574 243922 408642 243978
rect 408698 243922 408768 243978
rect 408448 243888 408768 243922
rect 439168 244350 439488 244384
rect 439168 244294 439238 244350
rect 439294 244294 439362 244350
rect 439418 244294 439488 244350
rect 439168 244226 439488 244294
rect 439168 244170 439238 244226
rect 439294 244170 439362 244226
rect 439418 244170 439488 244226
rect 439168 244102 439488 244170
rect 439168 244046 439238 244102
rect 439294 244046 439362 244102
rect 439418 244046 439488 244102
rect 439168 243978 439488 244046
rect 439168 243922 439238 243978
rect 439294 243922 439362 243978
rect 439418 243922 439488 243978
rect 439168 243888 439488 243922
rect 469888 244350 470208 244384
rect 469888 244294 469958 244350
rect 470014 244294 470082 244350
rect 470138 244294 470208 244350
rect 469888 244226 470208 244294
rect 469888 244170 469958 244226
rect 470014 244170 470082 244226
rect 470138 244170 470208 244226
rect 469888 244102 470208 244170
rect 469888 244046 469958 244102
rect 470014 244046 470082 244102
rect 470138 244046 470208 244102
rect 469888 243978 470208 244046
rect 469888 243922 469958 243978
rect 470014 243922 470082 243978
rect 470138 243922 470208 243978
rect 469888 243888 470208 243922
rect 500608 244350 500928 244384
rect 500608 244294 500678 244350
rect 500734 244294 500802 244350
rect 500858 244294 500928 244350
rect 500608 244226 500928 244294
rect 500608 244170 500678 244226
rect 500734 244170 500802 244226
rect 500858 244170 500928 244226
rect 500608 244102 500928 244170
rect 500608 244046 500678 244102
rect 500734 244046 500802 244102
rect 500858 244046 500928 244102
rect 500608 243978 500928 244046
rect 500608 243922 500678 243978
rect 500734 243922 500802 243978
rect 500858 243922 500928 243978
rect 500608 243888 500928 243922
rect 24448 238350 24768 238384
rect 24448 238294 24518 238350
rect 24574 238294 24642 238350
rect 24698 238294 24768 238350
rect 24448 238226 24768 238294
rect 24448 238170 24518 238226
rect 24574 238170 24642 238226
rect 24698 238170 24768 238226
rect 24448 238102 24768 238170
rect 24448 238046 24518 238102
rect 24574 238046 24642 238102
rect 24698 238046 24768 238102
rect 24448 237978 24768 238046
rect 24448 237922 24518 237978
rect 24574 237922 24642 237978
rect 24698 237922 24768 237978
rect 24448 237888 24768 237922
rect 55168 238350 55488 238384
rect 55168 238294 55238 238350
rect 55294 238294 55362 238350
rect 55418 238294 55488 238350
rect 55168 238226 55488 238294
rect 55168 238170 55238 238226
rect 55294 238170 55362 238226
rect 55418 238170 55488 238226
rect 55168 238102 55488 238170
rect 55168 238046 55238 238102
rect 55294 238046 55362 238102
rect 55418 238046 55488 238102
rect 55168 237978 55488 238046
rect 55168 237922 55238 237978
rect 55294 237922 55362 237978
rect 55418 237922 55488 237978
rect 55168 237888 55488 237922
rect 85888 238350 86208 238384
rect 85888 238294 85958 238350
rect 86014 238294 86082 238350
rect 86138 238294 86208 238350
rect 85888 238226 86208 238294
rect 85888 238170 85958 238226
rect 86014 238170 86082 238226
rect 86138 238170 86208 238226
rect 85888 238102 86208 238170
rect 85888 238046 85958 238102
rect 86014 238046 86082 238102
rect 86138 238046 86208 238102
rect 85888 237978 86208 238046
rect 85888 237922 85958 237978
rect 86014 237922 86082 237978
rect 86138 237922 86208 237978
rect 85888 237888 86208 237922
rect 116608 238350 116928 238384
rect 116608 238294 116678 238350
rect 116734 238294 116802 238350
rect 116858 238294 116928 238350
rect 116608 238226 116928 238294
rect 116608 238170 116678 238226
rect 116734 238170 116802 238226
rect 116858 238170 116928 238226
rect 116608 238102 116928 238170
rect 116608 238046 116678 238102
rect 116734 238046 116802 238102
rect 116858 238046 116928 238102
rect 116608 237978 116928 238046
rect 116608 237922 116678 237978
rect 116734 237922 116802 237978
rect 116858 237922 116928 237978
rect 116608 237888 116928 237922
rect 147328 238350 147648 238384
rect 147328 238294 147398 238350
rect 147454 238294 147522 238350
rect 147578 238294 147648 238350
rect 147328 238226 147648 238294
rect 147328 238170 147398 238226
rect 147454 238170 147522 238226
rect 147578 238170 147648 238226
rect 147328 238102 147648 238170
rect 147328 238046 147398 238102
rect 147454 238046 147522 238102
rect 147578 238046 147648 238102
rect 147328 237978 147648 238046
rect 147328 237922 147398 237978
rect 147454 237922 147522 237978
rect 147578 237922 147648 237978
rect 147328 237888 147648 237922
rect 178048 238350 178368 238384
rect 178048 238294 178118 238350
rect 178174 238294 178242 238350
rect 178298 238294 178368 238350
rect 178048 238226 178368 238294
rect 178048 238170 178118 238226
rect 178174 238170 178242 238226
rect 178298 238170 178368 238226
rect 178048 238102 178368 238170
rect 178048 238046 178118 238102
rect 178174 238046 178242 238102
rect 178298 238046 178368 238102
rect 178048 237978 178368 238046
rect 178048 237922 178118 237978
rect 178174 237922 178242 237978
rect 178298 237922 178368 237978
rect 178048 237888 178368 237922
rect 208768 238350 209088 238384
rect 208768 238294 208838 238350
rect 208894 238294 208962 238350
rect 209018 238294 209088 238350
rect 208768 238226 209088 238294
rect 208768 238170 208838 238226
rect 208894 238170 208962 238226
rect 209018 238170 209088 238226
rect 208768 238102 209088 238170
rect 208768 238046 208838 238102
rect 208894 238046 208962 238102
rect 209018 238046 209088 238102
rect 208768 237978 209088 238046
rect 208768 237922 208838 237978
rect 208894 237922 208962 237978
rect 209018 237922 209088 237978
rect 208768 237888 209088 237922
rect 239488 238350 239808 238384
rect 239488 238294 239558 238350
rect 239614 238294 239682 238350
rect 239738 238294 239808 238350
rect 239488 238226 239808 238294
rect 239488 238170 239558 238226
rect 239614 238170 239682 238226
rect 239738 238170 239808 238226
rect 239488 238102 239808 238170
rect 239488 238046 239558 238102
rect 239614 238046 239682 238102
rect 239738 238046 239808 238102
rect 239488 237978 239808 238046
rect 239488 237922 239558 237978
rect 239614 237922 239682 237978
rect 239738 237922 239808 237978
rect 239488 237888 239808 237922
rect 270208 238350 270528 238384
rect 270208 238294 270278 238350
rect 270334 238294 270402 238350
rect 270458 238294 270528 238350
rect 270208 238226 270528 238294
rect 270208 238170 270278 238226
rect 270334 238170 270402 238226
rect 270458 238170 270528 238226
rect 270208 238102 270528 238170
rect 270208 238046 270278 238102
rect 270334 238046 270402 238102
rect 270458 238046 270528 238102
rect 270208 237978 270528 238046
rect 270208 237922 270278 237978
rect 270334 237922 270402 237978
rect 270458 237922 270528 237978
rect 270208 237888 270528 237922
rect 300928 238350 301248 238384
rect 300928 238294 300998 238350
rect 301054 238294 301122 238350
rect 301178 238294 301248 238350
rect 300928 238226 301248 238294
rect 300928 238170 300998 238226
rect 301054 238170 301122 238226
rect 301178 238170 301248 238226
rect 300928 238102 301248 238170
rect 300928 238046 300998 238102
rect 301054 238046 301122 238102
rect 301178 238046 301248 238102
rect 300928 237978 301248 238046
rect 300928 237922 300998 237978
rect 301054 237922 301122 237978
rect 301178 237922 301248 237978
rect 300928 237888 301248 237922
rect 331648 238350 331968 238384
rect 331648 238294 331718 238350
rect 331774 238294 331842 238350
rect 331898 238294 331968 238350
rect 331648 238226 331968 238294
rect 331648 238170 331718 238226
rect 331774 238170 331842 238226
rect 331898 238170 331968 238226
rect 331648 238102 331968 238170
rect 331648 238046 331718 238102
rect 331774 238046 331842 238102
rect 331898 238046 331968 238102
rect 331648 237978 331968 238046
rect 331648 237922 331718 237978
rect 331774 237922 331842 237978
rect 331898 237922 331968 237978
rect 331648 237888 331968 237922
rect 362368 238350 362688 238384
rect 362368 238294 362438 238350
rect 362494 238294 362562 238350
rect 362618 238294 362688 238350
rect 362368 238226 362688 238294
rect 362368 238170 362438 238226
rect 362494 238170 362562 238226
rect 362618 238170 362688 238226
rect 362368 238102 362688 238170
rect 362368 238046 362438 238102
rect 362494 238046 362562 238102
rect 362618 238046 362688 238102
rect 362368 237978 362688 238046
rect 362368 237922 362438 237978
rect 362494 237922 362562 237978
rect 362618 237922 362688 237978
rect 362368 237888 362688 237922
rect 393088 238350 393408 238384
rect 393088 238294 393158 238350
rect 393214 238294 393282 238350
rect 393338 238294 393408 238350
rect 393088 238226 393408 238294
rect 393088 238170 393158 238226
rect 393214 238170 393282 238226
rect 393338 238170 393408 238226
rect 393088 238102 393408 238170
rect 393088 238046 393158 238102
rect 393214 238046 393282 238102
rect 393338 238046 393408 238102
rect 393088 237978 393408 238046
rect 393088 237922 393158 237978
rect 393214 237922 393282 237978
rect 393338 237922 393408 237978
rect 393088 237888 393408 237922
rect 423808 238350 424128 238384
rect 423808 238294 423878 238350
rect 423934 238294 424002 238350
rect 424058 238294 424128 238350
rect 423808 238226 424128 238294
rect 423808 238170 423878 238226
rect 423934 238170 424002 238226
rect 424058 238170 424128 238226
rect 423808 238102 424128 238170
rect 423808 238046 423878 238102
rect 423934 238046 424002 238102
rect 424058 238046 424128 238102
rect 423808 237978 424128 238046
rect 423808 237922 423878 237978
rect 423934 237922 424002 237978
rect 424058 237922 424128 237978
rect 423808 237888 424128 237922
rect 454528 238350 454848 238384
rect 454528 238294 454598 238350
rect 454654 238294 454722 238350
rect 454778 238294 454848 238350
rect 454528 238226 454848 238294
rect 454528 238170 454598 238226
rect 454654 238170 454722 238226
rect 454778 238170 454848 238226
rect 454528 238102 454848 238170
rect 454528 238046 454598 238102
rect 454654 238046 454722 238102
rect 454778 238046 454848 238102
rect 454528 237978 454848 238046
rect 454528 237922 454598 237978
rect 454654 237922 454722 237978
rect 454778 237922 454848 237978
rect 454528 237888 454848 237922
rect 485248 238350 485568 238384
rect 485248 238294 485318 238350
rect 485374 238294 485442 238350
rect 485498 238294 485568 238350
rect 485248 238226 485568 238294
rect 485248 238170 485318 238226
rect 485374 238170 485442 238226
rect 485498 238170 485568 238226
rect 485248 238102 485568 238170
rect 485248 238046 485318 238102
rect 485374 238046 485442 238102
rect 485498 238046 485568 238102
rect 485248 237978 485568 238046
rect 485248 237922 485318 237978
rect 485374 237922 485442 237978
rect 485498 237922 485568 237978
rect 485248 237888 485568 237922
rect 515968 238350 516288 238384
rect 515968 238294 516038 238350
rect 516094 238294 516162 238350
rect 516218 238294 516288 238350
rect 515968 238226 516288 238294
rect 515968 238170 516038 238226
rect 516094 238170 516162 238226
rect 516218 238170 516288 238226
rect 515968 238102 516288 238170
rect 515968 238046 516038 238102
rect 516094 238046 516162 238102
rect 516218 238046 516288 238102
rect 515968 237978 516288 238046
rect 515968 237922 516038 237978
rect 516094 237922 516162 237978
rect 516218 237922 516288 237978
rect 515968 237888 516288 237922
rect 525154 238350 525774 255922
rect 525154 238294 525250 238350
rect 525306 238294 525374 238350
rect 525430 238294 525498 238350
rect 525554 238294 525622 238350
rect 525678 238294 525774 238350
rect 525154 238226 525774 238294
rect 525154 238170 525250 238226
rect 525306 238170 525374 238226
rect 525430 238170 525498 238226
rect 525554 238170 525622 238226
rect 525678 238170 525774 238226
rect 525154 238102 525774 238170
rect 525154 238046 525250 238102
rect 525306 238046 525374 238102
rect 525430 238046 525498 238102
rect 525554 238046 525622 238102
rect 525678 238046 525774 238102
rect 525154 237978 525774 238046
rect 525154 237922 525250 237978
rect 525306 237922 525374 237978
rect 525430 237922 525498 237978
rect 525554 237922 525622 237978
rect 525678 237922 525774 237978
rect 6874 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 7494 226350
rect 6874 226226 7494 226294
rect 6874 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 7494 226226
rect 6874 226102 7494 226170
rect 6874 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 7494 226102
rect 6874 225978 7494 226046
rect 6874 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 7494 225978
rect 6874 208350 7494 225922
rect 39808 226350 40128 226384
rect 39808 226294 39878 226350
rect 39934 226294 40002 226350
rect 40058 226294 40128 226350
rect 39808 226226 40128 226294
rect 39808 226170 39878 226226
rect 39934 226170 40002 226226
rect 40058 226170 40128 226226
rect 39808 226102 40128 226170
rect 39808 226046 39878 226102
rect 39934 226046 40002 226102
rect 40058 226046 40128 226102
rect 39808 225978 40128 226046
rect 39808 225922 39878 225978
rect 39934 225922 40002 225978
rect 40058 225922 40128 225978
rect 39808 225888 40128 225922
rect 70528 226350 70848 226384
rect 70528 226294 70598 226350
rect 70654 226294 70722 226350
rect 70778 226294 70848 226350
rect 70528 226226 70848 226294
rect 70528 226170 70598 226226
rect 70654 226170 70722 226226
rect 70778 226170 70848 226226
rect 70528 226102 70848 226170
rect 70528 226046 70598 226102
rect 70654 226046 70722 226102
rect 70778 226046 70848 226102
rect 70528 225978 70848 226046
rect 70528 225922 70598 225978
rect 70654 225922 70722 225978
rect 70778 225922 70848 225978
rect 70528 225888 70848 225922
rect 101248 226350 101568 226384
rect 101248 226294 101318 226350
rect 101374 226294 101442 226350
rect 101498 226294 101568 226350
rect 101248 226226 101568 226294
rect 101248 226170 101318 226226
rect 101374 226170 101442 226226
rect 101498 226170 101568 226226
rect 101248 226102 101568 226170
rect 101248 226046 101318 226102
rect 101374 226046 101442 226102
rect 101498 226046 101568 226102
rect 101248 225978 101568 226046
rect 101248 225922 101318 225978
rect 101374 225922 101442 225978
rect 101498 225922 101568 225978
rect 101248 225888 101568 225922
rect 131968 226350 132288 226384
rect 131968 226294 132038 226350
rect 132094 226294 132162 226350
rect 132218 226294 132288 226350
rect 131968 226226 132288 226294
rect 131968 226170 132038 226226
rect 132094 226170 132162 226226
rect 132218 226170 132288 226226
rect 131968 226102 132288 226170
rect 131968 226046 132038 226102
rect 132094 226046 132162 226102
rect 132218 226046 132288 226102
rect 131968 225978 132288 226046
rect 131968 225922 132038 225978
rect 132094 225922 132162 225978
rect 132218 225922 132288 225978
rect 131968 225888 132288 225922
rect 162688 226350 163008 226384
rect 162688 226294 162758 226350
rect 162814 226294 162882 226350
rect 162938 226294 163008 226350
rect 162688 226226 163008 226294
rect 162688 226170 162758 226226
rect 162814 226170 162882 226226
rect 162938 226170 163008 226226
rect 162688 226102 163008 226170
rect 162688 226046 162758 226102
rect 162814 226046 162882 226102
rect 162938 226046 163008 226102
rect 162688 225978 163008 226046
rect 162688 225922 162758 225978
rect 162814 225922 162882 225978
rect 162938 225922 163008 225978
rect 162688 225888 163008 225922
rect 193408 226350 193728 226384
rect 193408 226294 193478 226350
rect 193534 226294 193602 226350
rect 193658 226294 193728 226350
rect 193408 226226 193728 226294
rect 193408 226170 193478 226226
rect 193534 226170 193602 226226
rect 193658 226170 193728 226226
rect 193408 226102 193728 226170
rect 193408 226046 193478 226102
rect 193534 226046 193602 226102
rect 193658 226046 193728 226102
rect 193408 225978 193728 226046
rect 193408 225922 193478 225978
rect 193534 225922 193602 225978
rect 193658 225922 193728 225978
rect 193408 225888 193728 225922
rect 224128 226350 224448 226384
rect 224128 226294 224198 226350
rect 224254 226294 224322 226350
rect 224378 226294 224448 226350
rect 224128 226226 224448 226294
rect 224128 226170 224198 226226
rect 224254 226170 224322 226226
rect 224378 226170 224448 226226
rect 224128 226102 224448 226170
rect 224128 226046 224198 226102
rect 224254 226046 224322 226102
rect 224378 226046 224448 226102
rect 224128 225978 224448 226046
rect 224128 225922 224198 225978
rect 224254 225922 224322 225978
rect 224378 225922 224448 225978
rect 224128 225888 224448 225922
rect 254848 226350 255168 226384
rect 254848 226294 254918 226350
rect 254974 226294 255042 226350
rect 255098 226294 255168 226350
rect 254848 226226 255168 226294
rect 254848 226170 254918 226226
rect 254974 226170 255042 226226
rect 255098 226170 255168 226226
rect 254848 226102 255168 226170
rect 254848 226046 254918 226102
rect 254974 226046 255042 226102
rect 255098 226046 255168 226102
rect 254848 225978 255168 226046
rect 254848 225922 254918 225978
rect 254974 225922 255042 225978
rect 255098 225922 255168 225978
rect 254848 225888 255168 225922
rect 285568 226350 285888 226384
rect 285568 226294 285638 226350
rect 285694 226294 285762 226350
rect 285818 226294 285888 226350
rect 285568 226226 285888 226294
rect 285568 226170 285638 226226
rect 285694 226170 285762 226226
rect 285818 226170 285888 226226
rect 285568 226102 285888 226170
rect 285568 226046 285638 226102
rect 285694 226046 285762 226102
rect 285818 226046 285888 226102
rect 285568 225978 285888 226046
rect 285568 225922 285638 225978
rect 285694 225922 285762 225978
rect 285818 225922 285888 225978
rect 285568 225888 285888 225922
rect 316288 226350 316608 226384
rect 316288 226294 316358 226350
rect 316414 226294 316482 226350
rect 316538 226294 316608 226350
rect 316288 226226 316608 226294
rect 316288 226170 316358 226226
rect 316414 226170 316482 226226
rect 316538 226170 316608 226226
rect 316288 226102 316608 226170
rect 316288 226046 316358 226102
rect 316414 226046 316482 226102
rect 316538 226046 316608 226102
rect 316288 225978 316608 226046
rect 316288 225922 316358 225978
rect 316414 225922 316482 225978
rect 316538 225922 316608 225978
rect 316288 225888 316608 225922
rect 347008 226350 347328 226384
rect 347008 226294 347078 226350
rect 347134 226294 347202 226350
rect 347258 226294 347328 226350
rect 347008 226226 347328 226294
rect 347008 226170 347078 226226
rect 347134 226170 347202 226226
rect 347258 226170 347328 226226
rect 347008 226102 347328 226170
rect 347008 226046 347078 226102
rect 347134 226046 347202 226102
rect 347258 226046 347328 226102
rect 347008 225978 347328 226046
rect 347008 225922 347078 225978
rect 347134 225922 347202 225978
rect 347258 225922 347328 225978
rect 347008 225888 347328 225922
rect 377728 226350 378048 226384
rect 377728 226294 377798 226350
rect 377854 226294 377922 226350
rect 377978 226294 378048 226350
rect 377728 226226 378048 226294
rect 377728 226170 377798 226226
rect 377854 226170 377922 226226
rect 377978 226170 378048 226226
rect 377728 226102 378048 226170
rect 377728 226046 377798 226102
rect 377854 226046 377922 226102
rect 377978 226046 378048 226102
rect 377728 225978 378048 226046
rect 377728 225922 377798 225978
rect 377854 225922 377922 225978
rect 377978 225922 378048 225978
rect 377728 225888 378048 225922
rect 408448 226350 408768 226384
rect 408448 226294 408518 226350
rect 408574 226294 408642 226350
rect 408698 226294 408768 226350
rect 408448 226226 408768 226294
rect 408448 226170 408518 226226
rect 408574 226170 408642 226226
rect 408698 226170 408768 226226
rect 408448 226102 408768 226170
rect 408448 226046 408518 226102
rect 408574 226046 408642 226102
rect 408698 226046 408768 226102
rect 408448 225978 408768 226046
rect 408448 225922 408518 225978
rect 408574 225922 408642 225978
rect 408698 225922 408768 225978
rect 408448 225888 408768 225922
rect 439168 226350 439488 226384
rect 439168 226294 439238 226350
rect 439294 226294 439362 226350
rect 439418 226294 439488 226350
rect 439168 226226 439488 226294
rect 439168 226170 439238 226226
rect 439294 226170 439362 226226
rect 439418 226170 439488 226226
rect 439168 226102 439488 226170
rect 439168 226046 439238 226102
rect 439294 226046 439362 226102
rect 439418 226046 439488 226102
rect 439168 225978 439488 226046
rect 439168 225922 439238 225978
rect 439294 225922 439362 225978
rect 439418 225922 439488 225978
rect 439168 225888 439488 225922
rect 469888 226350 470208 226384
rect 469888 226294 469958 226350
rect 470014 226294 470082 226350
rect 470138 226294 470208 226350
rect 469888 226226 470208 226294
rect 469888 226170 469958 226226
rect 470014 226170 470082 226226
rect 470138 226170 470208 226226
rect 469888 226102 470208 226170
rect 469888 226046 469958 226102
rect 470014 226046 470082 226102
rect 470138 226046 470208 226102
rect 469888 225978 470208 226046
rect 469888 225922 469958 225978
rect 470014 225922 470082 225978
rect 470138 225922 470208 225978
rect 469888 225888 470208 225922
rect 500608 226350 500928 226384
rect 500608 226294 500678 226350
rect 500734 226294 500802 226350
rect 500858 226294 500928 226350
rect 500608 226226 500928 226294
rect 500608 226170 500678 226226
rect 500734 226170 500802 226226
rect 500858 226170 500928 226226
rect 500608 226102 500928 226170
rect 500608 226046 500678 226102
rect 500734 226046 500802 226102
rect 500858 226046 500928 226102
rect 500608 225978 500928 226046
rect 500608 225922 500678 225978
rect 500734 225922 500802 225978
rect 500858 225922 500928 225978
rect 500608 225888 500928 225922
rect 24448 220350 24768 220384
rect 24448 220294 24518 220350
rect 24574 220294 24642 220350
rect 24698 220294 24768 220350
rect 24448 220226 24768 220294
rect 24448 220170 24518 220226
rect 24574 220170 24642 220226
rect 24698 220170 24768 220226
rect 24448 220102 24768 220170
rect 24448 220046 24518 220102
rect 24574 220046 24642 220102
rect 24698 220046 24768 220102
rect 24448 219978 24768 220046
rect 24448 219922 24518 219978
rect 24574 219922 24642 219978
rect 24698 219922 24768 219978
rect 24448 219888 24768 219922
rect 55168 220350 55488 220384
rect 55168 220294 55238 220350
rect 55294 220294 55362 220350
rect 55418 220294 55488 220350
rect 55168 220226 55488 220294
rect 55168 220170 55238 220226
rect 55294 220170 55362 220226
rect 55418 220170 55488 220226
rect 55168 220102 55488 220170
rect 55168 220046 55238 220102
rect 55294 220046 55362 220102
rect 55418 220046 55488 220102
rect 55168 219978 55488 220046
rect 55168 219922 55238 219978
rect 55294 219922 55362 219978
rect 55418 219922 55488 219978
rect 55168 219888 55488 219922
rect 85888 220350 86208 220384
rect 85888 220294 85958 220350
rect 86014 220294 86082 220350
rect 86138 220294 86208 220350
rect 85888 220226 86208 220294
rect 85888 220170 85958 220226
rect 86014 220170 86082 220226
rect 86138 220170 86208 220226
rect 85888 220102 86208 220170
rect 85888 220046 85958 220102
rect 86014 220046 86082 220102
rect 86138 220046 86208 220102
rect 85888 219978 86208 220046
rect 85888 219922 85958 219978
rect 86014 219922 86082 219978
rect 86138 219922 86208 219978
rect 85888 219888 86208 219922
rect 116608 220350 116928 220384
rect 116608 220294 116678 220350
rect 116734 220294 116802 220350
rect 116858 220294 116928 220350
rect 116608 220226 116928 220294
rect 116608 220170 116678 220226
rect 116734 220170 116802 220226
rect 116858 220170 116928 220226
rect 116608 220102 116928 220170
rect 116608 220046 116678 220102
rect 116734 220046 116802 220102
rect 116858 220046 116928 220102
rect 116608 219978 116928 220046
rect 116608 219922 116678 219978
rect 116734 219922 116802 219978
rect 116858 219922 116928 219978
rect 116608 219888 116928 219922
rect 147328 220350 147648 220384
rect 147328 220294 147398 220350
rect 147454 220294 147522 220350
rect 147578 220294 147648 220350
rect 147328 220226 147648 220294
rect 147328 220170 147398 220226
rect 147454 220170 147522 220226
rect 147578 220170 147648 220226
rect 147328 220102 147648 220170
rect 147328 220046 147398 220102
rect 147454 220046 147522 220102
rect 147578 220046 147648 220102
rect 147328 219978 147648 220046
rect 147328 219922 147398 219978
rect 147454 219922 147522 219978
rect 147578 219922 147648 219978
rect 147328 219888 147648 219922
rect 178048 220350 178368 220384
rect 178048 220294 178118 220350
rect 178174 220294 178242 220350
rect 178298 220294 178368 220350
rect 178048 220226 178368 220294
rect 178048 220170 178118 220226
rect 178174 220170 178242 220226
rect 178298 220170 178368 220226
rect 178048 220102 178368 220170
rect 178048 220046 178118 220102
rect 178174 220046 178242 220102
rect 178298 220046 178368 220102
rect 178048 219978 178368 220046
rect 178048 219922 178118 219978
rect 178174 219922 178242 219978
rect 178298 219922 178368 219978
rect 178048 219888 178368 219922
rect 208768 220350 209088 220384
rect 208768 220294 208838 220350
rect 208894 220294 208962 220350
rect 209018 220294 209088 220350
rect 208768 220226 209088 220294
rect 208768 220170 208838 220226
rect 208894 220170 208962 220226
rect 209018 220170 209088 220226
rect 208768 220102 209088 220170
rect 208768 220046 208838 220102
rect 208894 220046 208962 220102
rect 209018 220046 209088 220102
rect 208768 219978 209088 220046
rect 208768 219922 208838 219978
rect 208894 219922 208962 219978
rect 209018 219922 209088 219978
rect 208768 219888 209088 219922
rect 239488 220350 239808 220384
rect 239488 220294 239558 220350
rect 239614 220294 239682 220350
rect 239738 220294 239808 220350
rect 239488 220226 239808 220294
rect 239488 220170 239558 220226
rect 239614 220170 239682 220226
rect 239738 220170 239808 220226
rect 239488 220102 239808 220170
rect 239488 220046 239558 220102
rect 239614 220046 239682 220102
rect 239738 220046 239808 220102
rect 239488 219978 239808 220046
rect 239488 219922 239558 219978
rect 239614 219922 239682 219978
rect 239738 219922 239808 219978
rect 239488 219888 239808 219922
rect 270208 220350 270528 220384
rect 270208 220294 270278 220350
rect 270334 220294 270402 220350
rect 270458 220294 270528 220350
rect 270208 220226 270528 220294
rect 270208 220170 270278 220226
rect 270334 220170 270402 220226
rect 270458 220170 270528 220226
rect 270208 220102 270528 220170
rect 270208 220046 270278 220102
rect 270334 220046 270402 220102
rect 270458 220046 270528 220102
rect 270208 219978 270528 220046
rect 270208 219922 270278 219978
rect 270334 219922 270402 219978
rect 270458 219922 270528 219978
rect 270208 219888 270528 219922
rect 300928 220350 301248 220384
rect 300928 220294 300998 220350
rect 301054 220294 301122 220350
rect 301178 220294 301248 220350
rect 300928 220226 301248 220294
rect 300928 220170 300998 220226
rect 301054 220170 301122 220226
rect 301178 220170 301248 220226
rect 300928 220102 301248 220170
rect 300928 220046 300998 220102
rect 301054 220046 301122 220102
rect 301178 220046 301248 220102
rect 300928 219978 301248 220046
rect 300928 219922 300998 219978
rect 301054 219922 301122 219978
rect 301178 219922 301248 219978
rect 300928 219888 301248 219922
rect 331648 220350 331968 220384
rect 331648 220294 331718 220350
rect 331774 220294 331842 220350
rect 331898 220294 331968 220350
rect 331648 220226 331968 220294
rect 331648 220170 331718 220226
rect 331774 220170 331842 220226
rect 331898 220170 331968 220226
rect 331648 220102 331968 220170
rect 331648 220046 331718 220102
rect 331774 220046 331842 220102
rect 331898 220046 331968 220102
rect 331648 219978 331968 220046
rect 331648 219922 331718 219978
rect 331774 219922 331842 219978
rect 331898 219922 331968 219978
rect 331648 219888 331968 219922
rect 362368 220350 362688 220384
rect 362368 220294 362438 220350
rect 362494 220294 362562 220350
rect 362618 220294 362688 220350
rect 362368 220226 362688 220294
rect 362368 220170 362438 220226
rect 362494 220170 362562 220226
rect 362618 220170 362688 220226
rect 362368 220102 362688 220170
rect 362368 220046 362438 220102
rect 362494 220046 362562 220102
rect 362618 220046 362688 220102
rect 362368 219978 362688 220046
rect 362368 219922 362438 219978
rect 362494 219922 362562 219978
rect 362618 219922 362688 219978
rect 362368 219888 362688 219922
rect 393088 220350 393408 220384
rect 393088 220294 393158 220350
rect 393214 220294 393282 220350
rect 393338 220294 393408 220350
rect 393088 220226 393408 220294
rect 393088 220170 393158 220226
rect 393214 220170 393282 220226
rect 393338 220170 393408 220226
rect 393088 220102 393408 220170
rect 393088 220046 393158 220102
rect 393214 220046 393282 220102
rect 393338 220046 393408 220102
rect 393088 219978 393408 220046
rect 393088 219922 393158 219978
rect 393214 219922 393282 219978
rect 393338 219922 393408 219978
rect 393088 219888 393408 219922
rect 423808 220350 424128 220384
rect 423808 220294 423878 220350
rect 423934 220294 424002 220350
rect 424058 220294 424128 220350
rect 423808 220226 424128 220294
rect 423808 220170 423878 220226
rect 423934 220170 424002 220226
rect 424058 220170 424128 220226
rect 423808 220102 424128 220170
rect 423808 220046 423878 220102
rect 423934 220046 424002 220102
rect 424058 220046 424128 220102
rect 423808 219978 424128 220046
rect 423808 219922 423878 219978
rect 423934 219922 424002 219978
rect 424058 219922 424128 219978
rect 423808 219888 424128 219922
rect 454528 220350 454848 220384
rect 454528 220294 454598 220350
rect 454654 220294 454722 220350
rect 454778 220294 454848 220350
rect 454528 220226 454848 220294
rect 454528 220170 454598 220226
rect 454654 220170 454722 220226
rect 454778 220170 454848 220226
rect 454528 220102 454848 220170
rect 454528 220046 454598 220102
rect 454654 220046 454722 220102
rect 454778 220046 454848 220102
rect 454528 219978 454848 220046
rect 454528 219922 454598 219978
rect 454654 219922 454722 219978
rect 454778 219922 454848 219978
rect 454528 219888 454848 219922
rect 485248 220350 485568 220384
rect 485248 220294 485318 220350
rect 485374 220294 485442 220350
rect 485498 220294 485568 220350
rect 485248 220226 485568 220294
rect 485248 220170 485318 220226
rect 485374 220170 485442 220226
rect 485498 220170 485568 220226
rect 485248 220102 485568 220170
rect 485248 220046 485318 220102
rect 485374 220046 485442 220102
rect 485498 220046 485568 220102
rect 485248 219978 485568 220046
rect 485248 219922 485318 219978
rect 485374 219922 485442 219978
rect 485498 219922 485568 219978
rect 485248 219888 485568 219922
rect 515968 220350 516288 220384
rect 515968 220294 516038 220350
rect 516094 220294 516162 220350
rect 516218 220294 516288 220350
rect 515968 220226 516288 220294
rect 515968 220170 516038 220226
rect 516094 220170 516162 220226
rect 516218 220170 516288 220226
rect 515968 220102 516288 220170
rect 515968 220046 516038 220102
rect 516094 220046 516162 220102
rect 516218 220046 516288 220102
rect 515968 219978 516288 220046
rect 515968 219922 516038 219978
rect 516094 219922 516162 219978
rect 516218 219922 516288 219978
rect 515968 219888 516288 219922
rect 525154 220350 525774 237922
rect 525154 220294 525250 220350
rect 525306 220294 525374 220350
rect 525430 220294 525498 220350
rect 525554 220294 525622 220350
rect 525678 220294 525774 220350
rect 525154 220226 525774 220294
rect 525154 220170 525250 220226
rect 525306 220170 525374 220226
rect 525430 220170 525498 220226
rect 525554 220170 525622 220226
rect 525678 220170 525774 220226
rect 525154 220102 525774 220170
rect 525154 220046 525250 220102
rect 525306 220046 525374 220102
rect 525430 220046 525498 220102
rect 525554 220046 525622 220102
rect 525678 220046 525774 220102
rect 525154 219978 525774 220046
rect 525154 219922 525250 219978
rect 525306 219922 525374 219978
rect 525430 219922 525498 219978
rect 525554 219922 525622 219978
rect 525678 219922 525774 219978
rect 6874 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 7494 208350
rect 6874 208226 7494 208294
rect 6874 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 7494 208226
rect 6874 208102 7494 208170
rect 6874 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 7494 208102
rect 6874 207978 7494 208046
rect 6874 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 7494 207978
rect 6874 190350 7494 207922
rect 39808 208350 40128 208384
rect 39808 208294 39878 208350
rect 39934 208294 40002 208350
rect 40058 208294 40128 208350
rect 39808 208226 40128 208294
rect 39808 208170 39878 208226
rect 39934 208170 40002 208226
rect 40058 208170 40128 208226
rect 39808 208102 40128 208170
rect 39808 208046 39878 208102
rect 39934 208046 40002 208102
rect 40058 208046 40128 208102
rect 39808 207978 40128 208046
rect 39808 207922 39878 207978
rect 39934 207922 40002 207978
rect 40058 207922 40128 207978
rect 39808 207888 40128 207922
rect 70528 208350 70848 208384
rect 70528 208294 70598 208350
rect 70654 208294 70722 208350
rect 70778 208294 70848 208350
rect 70528 208226 70848 208294
rect 70528 208170 70598 208226
rect 70654 208170 70722 208226
rect 70778 208170 70848 208226
rect 70528 208102 70848 208170
rect 70528 208046 70598 208102
rect 70654 208046 70722 208102
rect 70778 208046 70848 208102
rect 70528 207978 70848 208046
rect 70528 207922 70598 207978
rect 70654 207922 70722 207978
rect 70778 207922 70848 207978
rect 70528 207888 70848 207922
rect 101248 208350 101568 208384
rect 101248 208294 101318 208350
rect 101374 208294 101442 208350
rect 101498 208294 101568 208350
rect 101248 208226 101568 208294
rect 101248 208170 101318 208226
rect 101374 208170 101442 208226
rect 101498 208170 101568 208226
rect 101248 208102 101568 208170
rect 101248 208046 101318 208102
rect 101374 208046 101442 208102
rect 101498 208046 101568 208102
rect 101248 207978 101568 208046
rect 101248 207922 101318 207978
rect 101374 207922 101442 207978
rect 101498 207922 101568 207978
rect 101248 207888 101568 207922
rect 131968 208350 132288 208384
rect 131968 208294 132038 208350
rect 132094 208294 132162 208350
rect 132218 208294 132288 208350
rect 131968 208226 132288 208294
rect 131968 208170 132038 208226
rect 132094 208170 132162 208226
rect 132218 208170 132288 208226
rect 131968 208102 132288 208170
rect 131968 208046 132038 208102
rect 132094 208046 132162 208102
rect 132218 208046 132288 208102
rect 131968 207978 132288 208046
rect 131968 207922 132038 207978
rect 132094 207922 132162 207978
rect 132218 207922 132288 207978
rect 131968 207888 132288 207922
rect 162688 208350 163008 208384
rect 162688 208294 162758 208350
rect 162814 208294 162882 208350
rect 162938 208294 163008 208350
rect 162688 208226 163008 208294
rect 162688 208170 162758 208226
rect 162814 208170 162882 208226
rect 162938 208170 163008 208226
rect 162688 208102 163008 208170
rect 162688 208046 162758 208102
rect 162814 208046 162882 208102
rect 162938 208046 163008 208102
rect 162688 207978 163008 208046
rect 162688 207922 162758 207978
rect 162814 207922 162882 207978
rect 162938 207922 163008 207978
rect 162688 207888 163008 207922
rect 193408 208350 193728 208384
rect 193408 208294 193478 208350
rect 193534 208294 193602 208350
rect 193658 208294 193728 208350
rect 193408 208226 193728 208294
rect 193408 208170 193478 208226
rect 193534 208170 193602 208226
rect 193658 208170 193728 208226
rect 193408 208102 193728 208170
rect 193408 208046 193478 208102
rect 193534 208046 193602 208102
rect 193658 208046 193728 208102
rect 193408 207978 193728 208046
rect 193408 207922 193478 207978
rect 193534 207922 193602 207978
rect 193658 207922 193728 207978
rect 193408 207888 193728 207922
rect 224128 208350 224448 208384
rect 224128 208294 224198 208350
rect 224254 208294 224322 208350
rect 224378 208294 224448 208350
rect 224128 208226 224448 208294
rect 224128 208170 224198 208226
rect 224254 208170 224322 208226
rect 224378 208170 224448 208226
rect 224128 208102 224448 208170
rect 224128 208046 224198 208102
rect 224254 208046 224322 208102
rect 224378 208046 224448 208102
rect 224128 207978 224448 208046
rect 224128 207922 224198 207978
rect 224254 207922 224322 207978
rect 224378 207922 224448 207978
rect 224128 207888 224448 207922
rect 254848 208350 255168 208384
rect 254848 208294 254918 208350
rect 254974 208294 255042 208350
rect 255098 208294 255168 208350
rect 254848 208226 255168 208294
rect 254848 208170 254918 208226
rect 254974 208170 255042 208226
rect 255098 208170 255168 208226
rect 254848 208102 255168 208170
rect 254848 208046 254918 208102
rect 254974 208046 255042 208102
rect 255098 208046 255168 208102
rect 254848 207978 255168 208046
rect 254848 207922 254918 207978
rect 254974 207922 255042 207978
rect 255098 207922 255168 207978
rect 254848 207888 255168 207922
rect 285568 208350 285888 208384
rect 285568 208294 285638 208350
rect 285694 208294 285762 208350
rect 285818 208294 285888 208350
rect 285568 208226 285888 208294
rect 285568 208170 285638 208226
rect 285694 208170 285762 208226
rect 285818 208170 285888 208226
rect 285568 208102 285888 208170
rect 285568 208046 285638 208102
rect 285694 208046 285762 208102
rect 285818 208046 285888 208102
rect 285568 207978 285888 208046
rect 285568 207922 285638 207978
rect 285694 207922 285762 207978
rect 285818 207922 285888 207978
rect 285568 207888 285888 207922
rect 316288 208350 316608 208384
rect 316288 208294 316358 208350
rect 316414 208294 316482 208350
rect 316538 208294 316608 208350
rect 316288 208226 316608 208294
rect 316288 208170 316358 208226
rect 316414 208170 316482 208226
rect 316538 208170 316608 208226
rect 316288 208102 316608 208170
rect 316288 208046 316358 208102
rect 316414 208046 316482 208102
rect 316538 208046 316608 208102
rect 316288 207978 316608 208046
rect 316288 207922 316358 207978
rect 316414 207922 316482 207978
rect 316538 207922 316608 207978
rect 316288 207888 316608 207922
rect 347008 208350 347328 208384
rect 347008 208294 347078 208350
rect 347134 208294 347202 208350
rect 347258 208294 347328 208350
rect 347008 208226 347328 208294
rect 347008 208170 347078 208226
rect 347134 208170 347202 208226
rect 347258 208170 347328 208226
rect 347008 208102 347328 208170
rect 347008 208046 347078 208102
rect 347134 208046 347202 208102
rect 347258 208046 347328 208102
rect 347008 207978 347328 208046
rect 347008 207922 347078 207978
rect 347134 207922 347202 207978
rect 347258 207922 347328 207978
rect 347008 207888 347328 207922
rect 377728 208350 378048 208384
rect 377728 208294 377798 208350
rect 377854 208294 377922 208350
rect 377978 208294 378048 208350
rect 377728 208226 378048 208294
rect 377728 208170 377798 208226
rect 377854 208170 377922 208226
rect 377978 208170 378048 208226
rect 377728 208102 378048 208170
rect 377728 208046 377798 208102
rect 377854 208046 377922 208102
rect 377978 208046 378048 208102
rect 377728 207978 378048 208046
rect 377728 207922 377798 207978
rect 377854 207922 377922 207978
rect 377978 207922 378048 207978
rect 377728 207888 378048 207922
rect 408448 208350 408768 208384
rect 408448 208294 408518 208350
rect 408574 208294 408642 208350
rect 408698 208294 408768 208350
rect 408448 208226 408768 208294
rect 408448 208170 408518 208226
rect 408574 208170 408642 208226
rect 408698 208170 408768 208226
rect 408448 208102 408768 208170
rect 408448 208046 408518 208102
rect 408574 208046 408642 208102
rect 408698 208046 408768 208102
rect 408448 207978 408768 208046
rect 408448 207922 408518 207978
rect 408574 207922 408642 207978
rect 408698 207922 408768 207978
rect 408448 207888 408768 207922
rect 439168 208350 439488 208384
rect 439168 208294 439238 208350
rect 439294 208294 439362 208350
rect 439418 208294 439488 208350
rect 439168 208226 439488 208294
rect 439168 208170 439238 208226
rect 439294 208170 439362 208226
rect 439418 208170 439488 208226
rect 439168 208102 439488 208170
rect 439168 208046 439238 208102
rect 439294 208046 439362 208102
rect 439418 208046 439488 208102
rect 439168 207978 439488 208046
rect 439168 207922 439238 207978
rect 439294 207922 439362 207978
rect 439418 207922 439488 207978
rect 439168 207888 439488 207922
rect 469888 208350 470208 208384
rect 469888 208294 469958 208350
rect 470014 208294 470082 208350
rect 470138 208294 470208 208350
rect 469888 208226 470208 208294
rect 469888 208170 469958 208226
rect 470014 208170 470082 208226
rect 470138 208170 470208 208226
rect 469888 208102 470208 208170
rect 469888 208046 469958 208102
rect 470014 208046 470082 208102
rect 470138 208046 470208 208102
rect 469888 207978 470208 208046
rect 469888 207922 469958 207978
rect 470014 207922 470082 207978
rect 470138 207922 470208 207978
rect 469888 207888 470208 207922
rect 500608 208350 500928 208384
rect 500608 208294 500678 208350
rect 500734 208294 500802 208350
rect 500858 208294 500928 208350
rect 500608 208226 500928 208294
rect 500608 208170 500678 208226
rect 500734 208170 500802 208226
rect 500858 208170 500928 208226
rect 500608 208102 500928 208170
rect 500608 208046 500678 208102
rect 500734 208046 500802 208102
rect 500858 208046 500928 208102
rect 500608 207978 500928 208046
rect 500608 207922 500678 207978
rect 500734 207922 500802 207978
rect 500858 207922 500928 207978
rect 500608 207888 500928 207922
rect 24448 202350 24768 202384
rect 24448 202294 24518 202350
rect 24574 202294 24642 202350
rect 24698 202294 24768 202350
rect 24448 202226 24768 202294
rect 24448 202170 24518 202226
rect 24574 202170 24642 202226
rect 24698 202170 24768 202226
rect 24448 202102 24768 202170
rect 24448 202046 24518 202102
rect 24574 202046 24642 202102
rect 24698 202046 24768 202102
rect 24448 201978 24768 202046
rect 24448 201922 24518 201978
rect 24574 201922 24642 201978
rect 24698 201922 24768 201978
rect 24448 201888 24768 201922
rect 55168 202350 55488 202384
rect 55168 202294 55238 202350
rect 55294 202294 55362 202350
rect 55418 202294 55488 202350
rect 55168 202226 55488 202294
rect 55168 202170 55238 202226
rect 55294 202170 55362 202226
rect 55418 202170 55488 202226
rect 55168 202102 55488 202170
rect 55168 202046 55238 202102
rect 55294 202046 55362 202102
rect 55418 202046 55488 202102
rect 55168 201978 55488 202046
rect 55168 201922 55238 201978
rect 55294 201922 55362 201978
rect 55418 201922 55488 201978
rect 55168 201888 55488 201922
rect 85888 202350 86208 202384
rect 85888 202294 85958 202350
rect 86014 202294 86082 202350
rect 86138 202294 86208 202350
rect 85888 202226 86208 202294
rect 85888 202170 85958 202226
rect 86014 202170 86082 202226
rect 86138 202170 86208 202226
rect 85888 202102 86208 202170
rect 85888 202046 85958 202102
rect 86014 202046 86082 202102
rect 86138 202046 86208 202102
rect 85888 201978 86208 202046
rect 85888 201922 85958 201978
rect 86014 201922 86082 201978
rect 86138 201922 86208 201978
rect 85888 201888 86208 201922
rect 116608 202350 116928 202384
rect 116608 202294 116678 202350
rect 116734 202294 116802 202350
rect 116858 202294 116928 202350
rect 116608 202226 116928 202294
rect 116608 202170 116678 202226
rect 116734 202170 116802 202226
rect 116858 202170 116928 202226
rect 116608 202102 116928 202170
rect 116608 202046 116678 202102
rect 116734 202046 116802 202102
rect 116858 202046 116928 202102
rect 116608 201978 116928 202046
rect 116608 201922 116678 201978
rect 116734 201922 116802 201978
rect 116858 201922 116928 201978
rect 116608 201888 116928 201922
rect 147328 202350 147648 202384
rect 147328 202294 147398 202350
rect 147454 202294 147522 202350
rect 147578 202294 147648 202350
rect 147328 202226 147648 202294
rect 147328 202170 147398 202226
rect 147454 202170 147522 202226
rect 147578 202170 147648 202226
rect 147328 202102 147648 202170
rect 147328 202046 147398 202102
rect 147454 202046 147522 202102
rect 147578 202046 147648 202102
rect 147328 201978 147648 202046
rect 147328 201922 147398 201978
rect 147454 201922 147522 201978
rect 147578 201922 147648 201978
rect 147328 201888 147648 201922
rect 178048 202350 178368 202384
rect 178048 202294 178118 202350
rect 178174 202294 178242 202350
rect 178298 202294 178368 202350
rect 178048 202226 178368 202294
rect 178048 202170 178118 202226
rect 178174 202170 178242 202226
rect 178298 202170 178368 202226
rect 178048 202102 178368 202170
rect 178048 202046 178118 202102
rect 178174 202046 178242 202102
rect 178298 202046 178368 202102
rect 178048 201978 178368 202046
rect 178048 201922 178118 201978
rect 178174 201922 178242 201978
rect 178298 201922 178368 201978
rect 178048 201888 178368 201922
rect 208768 202350 209088 202384
rect 208768 202294 208838 202350
rect 208894 202294 208962 202350
rect 209018 202294 209088 202350
rect 208768 202226 209088 202294
rect 208768 202170 208838 202226
rect 208894 202170 208962 202226
rect 209018 202170 209088 202226
rect 208768 202102 209088 202170
rect 208768 202046 208838 202102
rect 208894 202046 208962 202102
rect 209018 202046 209088 202102
rect 208768 201978 209088 202046
rect 208768 201922 208838 201978
rect 208894 201922 208962 201978
rect 209018 201922 209088 201978
rect 208768 201888 209088 201922
rect 239488 202350 239808 202384
rect 239488 202294 239558 202350
rect 239614 202294 239682 202350
rect 239738 202294 239808 202350
rect 239488 202226 239808 202294
rect 239488 202170 239558 202226
rect 239614 202170 239682 202226
rect 239738 202170 239808 202226
rect 239488 202102 239808 202170
rect 239488 202046 239558 202102
rect 239614 202046 239682 202102
rect 239738 202046 239808 202102
rect 239488 201978 239808 202046
rect 239488 201922 239558 201978
rect 239614 201922 239682 201978
rect 239738 201922 239808 201978
rect 239488 201888 239808 201922
rect 270208 202350 270528 202384
rect 270208 202294 270278 202350
rect 270334 202294 270402 202350
rect 270458 202294 270528 202350
rect 270208 202226 270528 202294
rect 270208 202170 270278 202226
rect 270334 202170 270402 202226
rect 270458 202170 270528 202226
rect 270208 202102 270528 202170
rect 270208 202046 270278 202102
rect 270334 202046 270402 202102
rect 270458 202046 270528 202102
rect 270208 201978 270528 202046
rect 270208 201922 270278 201978
rect 270334 201922 270402 201978
rect 270458 201922 270528 201978
rect 270208 201888 270528 201922
rect 300928 202350 301248 202384
rect 300928 202294 300998 202350
rect 301054 202294 301122 202350
rect 301178 202294 301248 202350
rect 300928 202226 301248 202294
rect 300928 202170 300998 202226
rect 301054 202170 301122 202226
rect 301178 202170 301248 202226
rect 300928 202102 301248 202170
rect 300928 202046 300998 202102
rect 301054 202046 301122 202102
rect 301178 202046 301248 202102
rect 300928 201978 301248 202046
rect 300928 201922 300998 201978
rect 301054 201922 301122 201978
rect 301178 201922 301248 201978
rect 300928 201888 301248 201922
rect 331648 202350 331968 202384
rect 331648 202294 331718 202350
rect 331774 202294 331842 202350
rect 331898 202294 331968 202350
rect 331648 202226 331968 202294
rect 331648 202170 331718 202226
rect 331774 202170 331842 202226
rect 331898 202170 331968 202226
rect 331648 202102 331968 202170
rect 331648 202046 331718 202102
rect 331774 202046 331842 202102
rect 331898 202046 331968 202102
rect 331648 201978 331968 202046
rect 331648 201922 331718 201978
rect 331774 201922 331842 201978
rect 331898 201922 331968 201978
rect 331648 201888 331968 201922
rect 362368 202350 362688 202384
rect 362368 202294 362438 202350
rect 362494 202294 362562 202350
rect 362618 202294 362688 202350
rect 362368 202226 362688 202294
rect 362368 202170 362438 202226
rect 362494 202170 362562 202226
rect 362618 202170 362688 202226
rect 362368 202102 362688 202170
rect 362368 202046 362438 202102
rect 362494 202046 362562 202102
rect 362618 202046 362688 202102
rect 362368 201978 362688 202046
rect 362368 201922 362438 201978
rect 362494 201922 362562 201978
rect 362618 201922 362688 201978
rect 362368 201888 362688 201922
rect 393088 202350 393408 202384
rect 393088 202294 393158 202350
rect 393214 202294 393282 202350
rect 393338 202294 393408 202350
rect 393088 202226 393408 202294
rect 393088 202170 393158 202226
rect 393214 202170 393282 202226
rect 393338 202170 393408 202226
rect 393088 202102 393408 202170
rect 393088 202046 393158 202102
rect 393214 202046 393282 202102
rect 393338 202046 393408 202102
rect 393088 201978 393408 202046
rect 393088 201922 393158 201978
rect 393214 201922 393282 201978
rect 393338 201922 393408 201978
rect 393088 201888 393408 201922
rect 423808 202350 424128 202384
rect 423808 202294 423878 202350
rect 423934 202294 424002 202350
rect 424058 202294 424128 202350
rect 423808 202226 424128 202294
rect 423808 202170 423878 202226
rect 423934 202170 424002 202226
rect 424058 202170 424128 202226
rect 423808 202102 424128 202170
rect 423808 202046 423878 202102
rect 423934 202046 424002 202102
rect 424058 202046 424128 202102
rect 423808 201978 424128 202046
rect 423808 201922 423878 201978
rect 423934 201922 424002 201978
rect 424058 201922 424128 201978
rect 423808 201888 424128 201922
rect 454528 202350 454848 202384
rect 454528 202294 454598 202350
rect 454654 202294 454722 202350
rect 454778 202294 454848 202350
rect 454528 202226 454848 202294
rect 454528 202170 454598 202226
rect 454654 202170 454722 202226
rect 454778 202170 454848 202226
rect 454528 202102 454848 202170
rect 454528 202046 454598 202102
rect 454654 202046 454722 202102
rect 454778 202046 454848 202102
rect 454528 201978 454848 202046
rect 454528 201922 454598 201978
rect 454654 201922 454722 201978
rect 454778 201922 454848 201978
rect 454528 201888 454848 201922
rect 485248 202350 485568 202384
rect 485248 202294 485318 202350
rect 485374 202294 485442 202350
rect 485498 202294 485568 202350
rect 485248 202226 485568 202294
rect 485248 202170 485318 202226
rect 485374 202170 485442 202226
rect 485498 202170 485568 202226
rect 485248 202102 485568 202170
rect 485248 202046 485318 202102
rect 485374 202046 485442 202102
rect 485498 202046 485568 202102
rect 485248 201978 485568 202046
rect 485248 201922 485318 201978
rect 485374 201922 485442 201978
rect 485498 201922 485568 201978
rect 485248 201888 485568 201922
rect 515968 202350 516288 202384
rect 515968 202294 516038 202350
rect 516094 202294 516162 202350
rect 516218 202294 516288 202350
rect 515968 202226 516288 202294
rect 515968 202170 516038 202226
rect 516094 202170 516162 202226
rect 516218 202170 516288 202226
rect 515968 202102 516288 202170
rect 515968 202046 516038 202102
rect 516094 202046 516162 202102
rect 516218 202046 516288 202102
rect 515968 201978 516288 202046
rect 515968 201922 516038 201978
rect 516094 201922 516162 201978
rect 516218 201922 516288 201978
rect 515968 201888 516288 201922
rect 525154 202350 525774 219922
rect 525154 202294 525250 202350
rect 525306 202294 525374 202350
rect 525430 202294 525498 202350
rect 525554 202294 525622 202350
rect 525678 202294 525774 202350
rect 525154 202226 525774 202294
rect 525154 202170 525250 202226
rect 525306 202170 525374 202226
rect 525430 202170 525498 202226
rect 525554 202170 525622 202226
rect 525678 202170 525774 202226
rect 525154 202102 525774 202170
rect 525154 202046 525250 202102
rect 525306 202046 525374 202102
rect 525430 202046 525498 202102
rect 525554 202046 525622 202102
rect 525678 202046 525774 202102
rect 525154 201978 525774 202046
rect 525154 201922 525250 201978
rect 525306 201922 525374 201978
rect 525430 201922 525498 201978
rect 525554 201922 525622 201978
rect 525678 201922 525774 201978
rect 6874 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 7494 190350
rect 6874 190226 7494 190294
rect 6874 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 7494 190226
rect 6874 190102 7494 190170
rect 6874 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 7494 190102
rect 6874 189978 7494 190046
rect 6874 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 7494 189978
rect 6874 172350 7494 189922
rect 39808 190350 40128 190384
rect 39808 190294 39878 190350
rect 39934 190294 40002 190350
rect 40058 190294 40128 190350
rect 39808 190226 40128 190294
rect 39808 190170 39878 190226
rect 39934 190170 40002 190226
rect 40058 190170 40128 190226
rect 39808 190102 40128 190170
rect 39808 190046 39878 190102
rect 39934 190046 40002 190102
rect 40058 190046 40128 190102
rect 39808 189978 40128 190046
rect 39808 189922 39878 189978
rect 39934 189922 40002 189978
rect 40058 189922 40128 189978
rect 39808 189888 40128 189922
rect 70528 190350 70848 190384
rect 70528 190294 70598 190350
rect 70654 190294 70722 190350
rect 70778 190294 70848 190350
rect 70528 190226 70848 190294
rect 70528 190170 70598 190226
rect 70654 190170 70722 190226
rect 70778 190170 70848 190226
rect 70528 190102 70848 190170
rect 70528 190046 70598 190102
rect 70654 190046 70722 190102
rect 70778 190046 70848 190102
rect 70528 189978 70848 190046
rect 70528 189922 70598 189978
rect 70654 189922 70722 189978
rect 70778 189922 70848 189978
rect 70528 189888 70848 189922
rect 101248 190350 101568 190384
rect 101248 190294 101318 190350
rect 101374 190294 101442 190350
rect 101498 190294 101568 190350
rect 101248 190226 101568 190294
rect 101248 190170 101318 190226
rect 101374 190170 101442 190226
rect 101498 190170 101568 190226
rect 101248 190102 101568 190170
rect 101248 190046 101318 190102
rect 101374 190046 101442 190102
rect 101498 190046 101568 190102
rect 101248 189978 101568 190046
rect 101248 189922 101318 189978
rect 101374 189922 101442 189978
rect 101498 189922 101568 189978
rect 101248 189888 101568 189922
rect 131968 190350 132288 190384
rect 131968 190294 132038 190350
rect 132094 190294 132162 190350
rect 132218 190294 132288 190350
rect 131968 190226 132288 190294
rect 131968 190170 132038 190226
rect 132094 190170 132162 190226
rect 132218 190170 132288 190226
rect 131968 190102 132288 190170
rect 131968 190046 132038 190102
rect 132094 190046 132162 190102
rect 132218 190046 132288 190102
rect 131968 189978 132288 190046
rect 131968 189922 132038 189978
rect 132094 189922 132162 189978
rect 132218 189922 132288 189978
rect 131968 189888 132288 189922
rect 162688 190350 163008 190384
rect 162688 190294 162758 190350
rect 162814 190294 162882 190350
rect 162938 190294 163008 190350
rect 162688 190226 163008 190294
rect 162688 190170 162758 190226
rect 162814 190170 162882 190226
rect 162938 190170 163008 190226
rect 162688 190102 163008 190170
rect 162688 190046 162758 190102
rect 162814 190046 162882 190102
rect 162938 190046 163008 190102
rect 162688 189978 163008 190046
rect 162688 189922 162758 189978
rect 162814 189922 162882 189978
rect 162938 189922 163008 189978
rect 162688 189888 163008 189922
rect 193408 190350 193728 190384
rect 193408 190294 193478 190350
rect 193534 190294 193602 190350
rect 193658 190294 193728 190350
rect 193408 190226 193728 190294
rect 193408 190170 193478 190226
rect 193534 190170 193602 190226
rect 193658 190170 193728 190226
rect 193408 190102 193728 190170
rect 193408 190046 193478 190102
rect 193534 190046 193602 190102
rect 193658 190046 193728 190102
rect 193408 189978 193728 190046
rect 193408 189922 193478 189978
rect 193534 189922 193602 189978
rect 193658 189922 193728 189978
rect 193408 189888 193728 189922
rect 224128 190350 224448 190384
rect 224128 190294 224198 190350
rect 224254 190294 224322 190350
rect 224378 190294 224448 190350
rect 224128 190226 224448 190294
rect 224128 190170 224198 190226
rect 224254 190170 224322 190226
rect 224378 190170 224448 190226
rect 224128 190102 224448 190170
rect 224128 190046 224198 190102
rect 224254 190046 224322 190102
rect 224378 190046 224448 190102
rect 224128 189978 224448 190046
rect 224128 189922 224198 189978
rect 224254 189922 224322 189978
rect 224378 189922 224448 189978
rect 224128 189888 224448 189922
rect 254848 190350 255168 190384
rect 254848 190294 254918 190350
rect 254974 190294 255042 190350
rect 255098 190294 255168 190350
rect 254848 190226 255168 190294
rect 254848 190170 254918 190226
rect 254974 190170 255042 190226
rect 255098 190170 255168 190226
rect 254848 190102 255168 190170
rect 254848 190046 254918 190102
rect 254974 190046 255042 190102
rect 255098 190046 255168 190102
rect 254848 189978 255168 190046
rect 254848 189922 254918 189978
rect 254974 189922 255042 189978
rect 255098 189922 255168 189978
rect 254848 189888 255168 189922
rect 285568 190350 285888 190384
rect 285568 190294 285638 190350
rect 285694 190294 285762 190350
rect 285818 190294 285888 190350
rect 285568 190226 285888 190294
rect 285568 190170 285638 190226
rect 285694 190170 285762 190226
rect 285818 190170 285888 190226
rect 285568 190102 285888 190170
rect 285568 190046 285638 190102
rect 285694 190046 285762 190102
rect 285818 190046 285888 190102
rect 285568 189978 285888 190046
rect 285568 189922 285638 189978
rect 285694 189922 285762 189978
rect 285818 189922 285888 189978
rect 285568 189888 285888 189922
rect 316288 190350 316608 190384
rect 316288 190294 316358 190350
rect 316414 190294 316482 190350
rect 316538 190294 316608 190350
rect 316288 190226 316608 190294
rect 316288 190170 316358 190226
rect 316414 190170 316482 190226
rect 316538 190170 316608 190226
rect 316288 190102 316608 190170
rect 316288 190046 316358 190102
rect 316414 190046 316482 190102
rect 316538 190046 316608 190102
rect 316288 189978 316608 190046
rect 316288 189922 316358 189978
rect 316414 189922 316482 189978
rect 316538 189922 316608 189978
rect 316288 189888 316608 189922
rect 347008 190350 347328 190384
rect 347008 190294 347078 190350
rect 347134 190294 347202 190350
rect 347258 190294 347328 190350
rect 347008 190226 347328 190294
rect 347008 190170 347078 190226
rect 347134 190170 347202 190226
rect 347258 190170 347328 190226
rect 347008 190102 347328 190170
rect 347008 190046 347078 190102
rect 347134 190046 347202 190102
rect 347258 190046 347328 190102
rect 347008 189978 347328 190046
rect 347008 189922 347078 189978
rect 347134 189922 347202 189978
rect 347258 189922 347328 189978
rect 347008 189888 347328 189922
rect 377728 190350 378048 190384
rect 377728 190294 377798 190350
rect 377854 190294 377922 190350
rect 377978 190294 378048 190350
rect 377728 190226 378048 190294
rect 377728 190170 377798 190226
rect 377854 190170 377922 190226
rect 377978 190170 378048 190226
rect 377728 190102 378048 190170
rect 377728 190046 377798 190102
rect 377854 190046 377922 190102
rect 377978 190046 378048 190102
rect 377728 189978 378048 190046
rect 377728 189922 377798 189978
rect 377854 189922 377922 189978
rect 377978 189922 378048 189978
rect 377728 189888 378048 189922
rect 408448 190350 408768 190384
rect 408448 190294 408518 190350
rect 408574 190294 408642 190350
rect 408698 190294 408768 190350
rect 408448 190226 408768 190294
rect 408448 190170 408518 190226
rect 408574 190170 408642 190226
rect 408698 190170 408768 190226
rect 408448 190102 408768 190170
rect 408448 190046 408518 190102
rect 408574 190046 408642 190102
rect 408698 190046 408768 190102
rect 408448 189978 408768 190046
rect 408448 189922 408518 189978
rect 408574 189922 408642 189978
rect 408698 189922 408768 189978
rect 408448 189888 408768 189922
rect 439168 190350 439488 190384
rect 439168 190294 439238 190350
rect 439294 190294 439362 190350
rect 439418 190294 439488 190350
rect 439168 190226 439488 190294
rect 439168 190170 439238 190226
rect 439294 190170 439362 190226
rect 439418 190170 439488 190226
rect 439168 190102 439488 190170
rect 439168 190046 439238 190102
rect 439294 190046 439362 190102
rect 439418 190046 439488 190102
rect 439168 189978 439488 190046
rect 439168 189922 439238 189978
rect 439294 189922 439362 189978
rect 439418 189922 439488 189978
rect 439168 189888 439488 189922
rect 469888 190350 470208 190384
rect 469888 190294 469958 190350
rect 470014 190294 470082 190350
rect 470138 190294 470208 190350
rect 469888 190226 470208 190294
rect 469888 190170 469958 190226
rect 470014 190170 470082 190226
rect 470138 190170 470208 190226
rect 469888 190102 470208 190170
rect 469888 190046 469958 190102
rect 470014 190046 470082 190102
rect 470138 190046 470208 190102
rect 469888 189978 470208 190046
rect 469888 189922 469958 189978
rect 470014 189922 470082 189978
rect 470138 189922 470208 189978
rect 469888 189888 470208 189922
rect 500608 190350 500928 190384
rect 500608 190294 500678 190350
rect 500734 190294 500802 190350
rect 500858 190294 500928 190350
rect 500608 190226 500928 190294
rect 500608 190170 500678 190226
rect 500734 190170 500802 190226
rect 500858 190170 500928 190226
rect 500608 190102 500928 190170
rect 500608 190046 500678 190102
rect 500734 190046 500802 190102
rect 500858 190046 500928 190102
rect 500608 189978 500928 190046
rect 500608 189922 500678 189978
rect 500734 189922 500802 189978
rect 500858 189922 500928 189978
rect 500608 189888 500928 189922
rect 24448 184350 24768 184384
rect 24448 184294 24518 184350
rect 24574 184294 24642 184350
rect 24698 184294 24768 184350
rect 24448 184226 24768 184294
rect 24448 184170 24518 184226
rect 24574 184170 24642 184226
rect 24698 184170 24768 184226
rect 24448 184102 24768 184170
rect 24448 184046 24518 184102
rect 24574 184046 24642 184102
rect 24698 184046 24768 184102
rect 24448 183978 24768 184046
rect 24448 183922 24518 183978
rect 24574 183922 24642 183978
rect 24698 183922 24768 183978
rect 24448 183888 24768 183922
rect 55168 184350 55488 184384
rect 55168 184294 55238 184350
rect 55294 184294 55362 184350
rect 55418 184294 55488 184350
rect 55168 184226 55488 184294
rect 55168 184170 55238 184226
rect 55294 184170 55362 184226
rect 55418 184170 55488 184226
rect 55168 184102 55488 184170
rect 55168 184046 55238 184102
rect 55294 184046 55362 184102
rect 55418 184046 55488 184102
rect 55168 183978 55488 184046
rect 55168 183922 55238 183978
rect 55294 183922 55362 183978
rect 55418 183922 55488 183978
rect 55168 183888 55488 183922
rect 85888 184350 86208 184384
rect 85888 184294 85958 184350
rect 86014 184294 86082 184350
rect 86138 184294 86208 184350
rect 85888 184226 86208 184294
rect 85888 184170 85958 184226
rect 86014 184170 86082 184226
rect 86138 184170 86208 184226
rect 85888 184102 86208 184170
rect 85888 184046 85958 184102
rect 86014 184046 86082 184102
rect 86138 184046 86208 184102
rect 85888 183978 86208 184046
rect 85888 183922 85958 183978
rect 86014 183922 86082 183978
rect 86138 183922 86208 183978
rect 85888 183888 86208 183922
rect 116608 184350 116928 184384
rect 116608 184294 116678 184350
rect 116734 184294 116802 184350
rect 116858 184294 116928 184350
rect 116608 184226 116928 184294
rect 116608 184170 116678 184226
rect 116734 184170 116802 184226
rect 116858 184170 116928 184226
rect 116608 184102 116928 184170
rect 116608 184046 116678 184102
rect 116734 184046 116802 184102
rect 116858 184046 116928 184102
rect 116608 183978 116928 184046
rect 116608 183922 116678 183978
rect 116734 183922 116802 183978
rect 116858 183922 116928 183978
rect 116608 183888 116928 183922
rect 147328 184350 147648 184384
rect 147328 184294 147398 184350
rect 147454 184294 147522 184350
rect 147578 184294 147648 184350
rect 147328 184226 147648 184294
rect 147328 184170 147398 184226
rect 147454 184170 147522 184226
rect 147578 184170 147648 184226
rect 147328 184102 147648 184170
rect 147328 184046 147398 184102
rect 147454 184046 147522 184102
rect 147578 184046 147648 184102
rect 147328 183978 147648 184046
rect 147328 183922 147398 183978
rect 147454 183922 147522 183978
rect 147578 183922 147648 183978
rect 147328 183888 147648 183922
rect 178048 184350 178368 184384
rect 178048 184294 178118 184350
rect 178174 184294 178242 184350
rect 178298 184294 178368 184350
rect 178048 184226 178368 184294
rect 178048 184170 178118 184226
rect 178174 184170 178242 184226
rect 178298 184170 178368 184226
rect 178048 184102 178368 184170
rect 178048 184046 178118 184102
rect 178174 184046 178242 184102
rect 178298 184046 178368 184102
rect 178048 183978 178368 184046
rect 178048 183922 178118 183978
rect 178174 183922 178242 183978
rect 178298 183922 178368 183978
rect 178048 183888 178368 183922
rect 208768 184350 209088 184384
rect 208768 184294 208838 184350
rect 208894 184294 208962 184350
rect 209018 184294 209088 184350
rect 208768 184226 209088 184294
rect 208768 184170 208838 184226
rect 208894 184170 208962 184226
rect 209018 184170 209088 184226
rect 208768 184102 209088 184170
rect 208768 184046 208838 184102
rect 208894 184046 208962 184102
rect 209018 184046 209088 184102
rect 208768 183978 209088 184046
rect 208768 183922 208838 183978
rect 208894 183922 208962 183978
rect 209018 183922 209088 183978
rect 208768 183888 209088 183922
rect 239488 184350 239808 184384
rect 239488 184294 239558 184350
rect 239614 184294 239682 184350
rect 239738 184294 239808 184350
rect 239488 184226 239808 184294
rect 239488 184170 239558 184226
rect 239614 184170 239682 184226
rect 239738 184170 239808 184226
rect 239488 184102 239808 184170
rect 239488 184046 239558 184102
rect 239614 184046 239682 184102
rect 239738 184046 239808 184102
rect 239488 183978 239808 184046
rect 239488 183922 239558 183978
rect 239614 183922 239682 183978
rect 239738 183922 239808 183978
rect 239488 183888 239808 183922
rect 270208 184350 270528 184384
rect 270208 184294 270278 184350
rect 270334 184294 270402 184350
rect 270458 184294 270528 184350
rect 270208 184226 270528 184294
rect 270208 184170 270278 184226
rect 270334 184170 270402 184226
rect 270458 184170 270528 184226
rect 270208 184102 270528 184170
rect 270208 184046 270278 184102
rect 270334 184046 270402 184102
rect 270458 184046 270528 184102
rect 270208 183978 270528 184046
rect 270208 183922 270278 183978
rect 270334 183922 270402 183978
rect 270458 183922 270528 183978
rect 270208 183888 270528 183922
rect 300928 184350 301248 184384
rect 300928 184294 300998 184350
rect 301054 184294 301122 184350
rect 301178 184294 301248 184350
rect 300928 184226 301248 184294
rect 300928 184170 300998 184226
rect 301054 184170 301122 184226
rect 301178 184170 301248 184226
rect 300928 184102 301248 184170
rect 300928 184046 300998 184102
rect 301054 184046 301122 184102
rect 301178 184046 301248 184102
rect 300928 183978 301248 184046
rect 300928 183922 300998 183978
rect 301054 183922 301122 183978
rect 301178 183922 301248 183978
rect 300928 183888 301248 183922
rect 331648 184350 331968 184384
rect 331648 184294 331718 184350
rect 331774 184294 331842 184350
rect 331898 184294 331968 184350
rect 331648 184226 331968 184294
rect 331648 184170 331718 184226
rect 331774 184170 331842 184226
rect 331898 184170 331968 184226
rect 331648 184102 331968 184170
rect 331648 184046 331718 184102
rect 331774 184046 331842 184102
rect 331898 184046 331968 184102
rect 331648 183978 331968 184046
rect 331648 183922 331718 183978
rect 331774 183922 331842 183978
rect 331898 183922 331968 183978
rect 331648 183888 331968 183922
rect 362368 184350 362688 184384
rect 362368 184294 362438 184350
rect 362494 184294 362562 184350
rect 362618 184294 362688 184350
rect 362368 184226 362688 184294
rect 362368 184170 362438 184226
rect 362494 184170 362562 184226
rect 362618 184170 362688 184226
rect 362368 184102 362688 184170
rect 362368 184046 362438 184102
rect 362494 184046 362562 184102
rect 362618 184046 362688 184102
rect 362368 183978 362688 184046
rect 362368 183922 362438 183978
rect 362494 183922 362562 183978
rect 362618 183922 362688 183978
rect 362368 183888 362688 183922
rect 393088 184350 393408 184384
rect 393088 184294 393158 184350
rect 393214 184294 393282 184350
rect 393338 184294 393408 184350
rect 393088 184226 393408 184294
rect 393088 184170 393158 184226
rect 393214 184170 393282 184226
rect 393338 184170 393408 184226
rect 393088 184102 393408 184170
rect 393088 184046 393158 184102
rect 393214 184046 393282 184102
rect 393338 184046 393408 184102
rect 393088 183978 393408 184046
rect 393088 183922 393158 183978
rect 393214 183922 393282 183978
rect 393338 183922 393408 183978
rect 393088 183888 393408 183922
rect 423808 184350 424128 184384
rect 423808 184294 423878 184350
rect 423934 184294 424002 184350
rect 424058 184294 424128 184350
rect 423808 184226 424128 184294
rect 423808 184170 423878 184226
rect 423934 184170 424002 184226
rect 424058 184170 424128 184226
rect 423808 184102 424128 184170
rect 423808 184046 423878 184102
rect 423934 184046 424002 184102
rect 424058 184046 424128 184102
rect 423808 183978 424128 184046
rect 423808 183922 423878 183978
rect 423934 183922 424002 183978
rect 424058 183922 424128 183978
rect 423808 183888 424128 183922
rect 454528 184350 454848 184384
rect 454528 184294 454598 184350
rect 454654 184294 454722 184350
rect 454778 184294 454848 184350
rect 454528 184226 454848 184294
rect 454528 184170 454598 184226
rect 454654 184170 454722 184226
rect 454778 184170 454848 184226
rect 454528 184102 454848 184170
rect 454528 184046 454598 184102
rect 454654 184046 454722 184102
rect 454778 184046 454848 184102
rect 454528 183978 454848 184046
rect 454528 183922 454598 183978
rect 454654 183922 454722 183978
rect 454778 183922 454848 183978
rect 454528 183888 454848 183922
rect 485248 184350 485568 184384
rect 485248 184294 485318 184350
rect 485374 184294 485442 184350
rect 485498 184294 485568 184350
rect 485248 184226 485568 184294
rect 485248 184170 485318 184226
rect 485374 184170 485442 184226
rect 485498 184170 485568 184226
rect 485248 184102 485568 184170
rect 485248 184046 485318 184102
rect 485374 184046 485442 184102
rect 485498 184046 485568 184102
rect 485248 183978 485568 184046
rect 485248 183922 485318 183978
rect 485374 183922 485442 183978
rect 485498 183922 485568 183978
rect 485248 183888 485568 183922
rect 515968 184350 516288 184384
rect 515968 184294 516038 184350
rect 516094 184294 516162 184350
rect 516218 184294 516288 184350
rect 515968 184226 516288 184294
rect 515968 184170 516038 184226
rect 516094 184170 516162 184226
rect 516218 184170 516288 184226
rect 515968 184102 516288 184170
rect 515968 184046 516038 184102
rect 516094 184046 516162 184102
rect 516218 184046 516288 184102
rect 515968 183978 516288 184046
rect 515968 183922 516038 183978
rect 516094 183922 516162 183978
rect 516218 183922 516288 183978
rect 515968 183888 516288 183922
rect 525154 184350 525774 201922
rect 525154 184294 525250 184350
rect 525306 184294 525374 184350
rect 525430 184294 525498 184350
rect 525554 184294 525622 184350
rect 525678 184294 525774 184350
rect 525154 184226 525774 184294
rect 525154 184170 525250 184226
rect 525306 184170 525374 184226
rect 525430 184170 525498 184226
rect 525554 184170 525622 184226
rect 525678 184170 525774 184226
rect 525154 184102 525774 184170
rect 525154 184046 525250 184102
rect 525306 184046 525374 184102
rect 525430 184046 525498 184102
rect 525554 184046 525622 184102
rect 525678 184046 525774 184102
rect 525154 183978 525774 184046
rect 525154 183922 525250 183978
rect 525306 183922 525374 183978
rect 525430 183922 525498 183978
rect 525554 183922 525622 183978
rect 525678 183922 525774 183978
rect 6874 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 7494 172350
rect 6874 172226 7494 172294
rect 6874 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 7494 172226
rect 6874 172102 7494 172170
rect 6874 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 7494 172102
rect 6874 171978 7494 172046
rect 6874 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 7494 171978
rect 6874 154350 7494 171922
rect 39808 172350 40128 172384
rect 39808 172294 39878 172350
rect 39934 172294 40002 172350
rect 40058 172294 40128 172350
rect 39808 172226 40128 172294
rect 39808 172170 39878 172226
rect 39934 172170 40002 172226
rect 40058 172170 40128 172226
rect 39808 172102 40128 172170
rect 39808 172046 39878 172102
rect 39934 172046 40002 172102
rect 40058 172046 40128 172102
rect 39808 171978 40128 172046
rect 39808 171922 39878 171978
rect 39934 171922 40002 171978
rect 40058 171922 40128 171978
rect 39808 171888 40128 171922
rect 70528 172350 70848 172384
rect 70528 172294 70598 172350
rect 70654 172294 70722 172350
rect 70778 172294 70848 172350
rect 70528 172226 70848 172294
rect 70528 172170 70598 172226
rect 70654 172170 70722 172226
rect 70778 172170 70848 172226
rect 70528 172102 70848 172170
rect 70528 172046 70598 172102
rect 70654 172046 70722 172102
rect 70778 172046 70848 172102
rect 70528 171978 70848 172046
rect 70528 171922 70598 171978
rect 70654 171922 70722 171978
rect 70778 171922 70848 171978
rect 70528 171888 70848 171922
rect 101248 172350 101568 172384
rect 101248 172294 101318 172350
rect 101374 172294 101442 172350
rect 101498 172294 101568 172350
rect 101248 172226 101568 172294
rect 101248 172170 101318 172226
rect 101374 172170 101442 172226
rect 101498 172170 101568 172226
rect 101248 172102 101568 172170
rect 101248 172046 101318 172102
rect 101374 172046 101442 172102
rect 101498 172046 101568 172102
rect 101248 171978 101568 172046
rect 101248 171922 101318 171978
rect 101374 171922 101442 171978
rect 101498 171922 101568 171978
rect 101248 171888 101568 171922
rect 131968 172350 132288 172384
rect 131968 172294 132038 172350
rect 132094 172294 132162 172350
rect 132218 172294 132288 172350
rect 131968 172226 132288 172294
rect 131968 172170 132038 172226
rect 132094 172170 132162 172226
rect 132218 172170 132288 172226
rect 131968 172102 132288 172170
rect 131968 172046 132038 172102
rect 132094 172046 132162 172102
rect 132218 172046 132288 172102
rect 131968 171978 132288 172046
rect 131968 171922 132038 171978
rect 132094 171922 132162 171978
rect 132218 171922 132288 171978
rect 131968 171888 132288 171922
rect 162688 172350 163008 172384
rect 162688 172294 162758 172350
rect 162814 172294 162882 172350
rect 162938 172294 163008 172350
rect 162688 172226 163008 172294
rect 162688 172170 162758 172226
rect 162814 172170 162882 172226
rect 162938 172170 163008 172226
rect 162688 172102 163008 172170
rect 162688 172046 162758 172102
rect 162814 172046 162882 172102
rect 162938 172046 163008 172102
rect 162688 171978 163008 172046
rect 162688 171922 162758 171978
rect 162814 171922 162882 171978
rect 162938 171922 163008 171978
rect 162688 171888 163008 171922
rect 193408 172350 193728 172384
rect 193408 172294 193478 172350
rect 193534 172294 193602 172350
rect 193658 172294 193728 172350
rect 193408 172226 193728 172294
rect 193408 172170 193478 172226
rect 193534 172170 193602 172226
rect 193658 172170 193728 172226
rect 193408 172102 193728 172170
rect 193408 172046 193478 172102
rect 193534 172046 193602 172102
rect 193658 172046 193728 172102
rect 193408 171978 193728 172046
rect 193408 171922 193478 171978
rect 193534 171922 193602 171978
rect 193658 171922 193728 171978
rect 193408 171888 193728 171922
rect 224128 172350 224448 172384
rect 224128 172294 224198 172350
rect 224254 172294 224322 172350
rect 224378 172294 224448 172350
rect 224128 172226 224448 172294
rect 224128 172170 224198 172226
rect 224254 172170 224322 172226
rect 224378 172170 224448 172226
rect 224128 172102 224448 172170
rect 224128 172046 224198 172102
rect 224254 172046 224322 172102
rect 224378 172046 224448 172102
rect 224128 171978 224448 172046
rect 224128 171922 224198 171978
rect 224254 171922 224322 171978
rect 224378 171922 224448 171978
rect 224128 171888 224448 171922
rect 254848 172350 255168 172384
rect 254848 172294 254918 172350
rect 254974 172294 255042 172350
rect 255098 172294 255168 172350
rect 254848 172226 255168 172294
rect 254848 172170 254918 172226
rect 254974 172170 255042 172226
rect 255098 172170 255168 172226
rect 254848 172102 255168 172170
rect 254848 172046 254918 172102
rect 254974 172046 255042 172102
rect 255098 172046 255168 172102
rect 254848 171978 255168 172046
rect 254848 171922 254918 171978
rect 254974 171922 255042 171978
rect 255098 171922 255168 171978
rect 254848 171888 255168 171922
rect 285568 172350 285888 172384
rect 285568 172294 285638 172350
rect 285694 172294 285762 172350
rect 285818 172294 285888 172350
rect 285568 172226 285888 172294
rect 285568 172170 285638 172226
rect 285694 172170 285762 172226
rect 285818 172170 285888 172226
rect 285568 172102 285888 172170
rect 285568 172046 285638 172102
rect 285694 172046 285762 172102
rect 285818 172046 285888 172102
rect 285568 171978 285888 172046
rect 285568 171922 285638 171978
rect 285694 171922 285762 171978
rect 285818 171922 285888 171978
rect 285568 171888 285888 171922
rect 316288 172350 316608 172384
rect 316288 172294 316358 172350
rect 316414 172294 316482 172350
rect 316538 172294 316608 172350
rect 316288 172226 316608 172294
rect 316288 172170 316358 172226
rect 316414 172170 316482 172226
rect 316538 172170 316608 172226
rect 316288 172102 316608 172170
rect 316288 172046 316358 172102
rect 316414 172046 316482 172102
rect 316538 172046 316608 172102
rect 316288 171978 316608 172046
rect 316288 171922 316358 171978
rect 316414 171922 316482 171978
rect 316538 171922 316608 171978
rect 316288 171888 316608 171922
rect 347008 172350 347328 172384
rect 347008 172294 347078 172350
rect 347134 172294 347202 172350
rect 347258 172294 347328 172350
rect 347008 172226 347328 172294
rect 347008 172170 347078 172226
rect 347134 172170 347202 172226
rect 347258 172170 347328 172226
rect 347008 172102 347328 172170
rect 347008 172046 347078 172102
rect 347134 172046 347202 172102
rect 347258 172046 347328 172102
rect 347008 171978 347328 172046
rect 347008 171922 347078 171978
rect 347134 171922 347202 171978
rect 347258 171922 347328 171978
rect 347008 171888 347328 171922
rect 377728 172350 378048 172384
rect 377728 172294 377798 172350
rect 377854 172294 377922 172350
rect 377978 172294 378048 172350
rect 377728 172226 378048 172294
rect 377728 172170 377798 172226
rect 377854 172170 377922 172226
rect 377978 172170 378048 172226
rect 377728 172102 378048 172170
rect 377728 172046 377798 172102
rect 377854 172046 377922 172102
rect 377978 172046 378048 172102
rect 377728 171978 378048 172046
rect 377728 171922 377798 171978
rect 377854 171922 377922 171978
rect 377978 171922 378048 171978
rect 377728 171888 378048 171922
rect 408448 172350 408768 172384
rect 408448 172294 408518 172350
rect 408574 172294 408642 172350
rect 408698 172294 408768 172350
rect 408448 172226 408768 172294
rect 408448 172170 408518 172226
rect 408574 172170 408642 172226
rect 408698 172170 408768 172226
rect 408448 172102 408768 172170
rect 408448 172046 408518 172102
rect 408574 172046 408642 172102
rect 408698 172046 408768 172102
rect 408448 171978 408768 172046
rect 408448 171922 408518 171978
rect 408574 171922 408642 171978
rect 408698 171922 408768 171978
rect 408448 171888 408768 171922
rect 439168 172350 439488 172384
rect 439168 172294 439238 172350
rect 439294 172294 439362 172350
rect 439418 172294 439488 172350
rect 439168 172226 439488 172294
rect 439168 172170 439238 172226
rect 439294 172170 439362 172226
rect 439418 172170 439488 172226
rect 439168 172102 439488 172170
rect 439168 172046 439238 172102
rect 439294 172046 439362 172102
rect 439418 172046 439488 172102
rect 439168 171978 439488 172046
rect 439168 171922 439238 171978
rect 439294 171922 439362 171978
rect 439418 171922 439488 171978
rect 439168 171888 439488 171922
rect 469888 172350 470208 172384
rect 469888 172294 469958 172350
rect 470014 172294 470082 172350
rect 470138 172294 470208 172350
rect 469888 172226 470208 172294
rect 469888 172170 469958 172226
rect 470014 172170 470082 172226
rect 470138 172170 470208 172226
rect 469888 172102 470208 172170
rect 469888 172046 469958 172102
rect 470014 172046 470082 172102
rect 470138 172046 470208 172102
rect 469888 171978 470208 172046
rect 469888 171922 469958 171978
rect 470014 171922 470082 171978
rect 470138 171922 470208 171978
rect 469888 171888 470208 171922
rect 500608 172350 500928 172384
rect 500608 172294 500678 172350
rect 500734 172294 500802 172350
rect 500858 172294 500928 172350
rect 500608 172226 500928 172294
rect 500608 172170 500678 172226
rect 500734 172170 500802 172226
rect 500858 172170 500928 172226
rect 500608 172102 500928 172170
rect 500608 172046 500678 172102
rect 500734 172046 500802 172102
rect 500858 172046 500928 172102
rect 500608 171978 500928 172046
rect 500608 171922 500678 171978
rect 500734 171922 500802 171978
rect 500858 171922 500928 171978
rect 500608 171888 500928 171922
rect 24448 166350 24768 166384
rect 24448 166294 24518 166350
rect 24574 166294 24642 166350
rect 24698 166294 24768 166350
rect 24448 166226 24768 166294
rect 24448 166170 24518 166226
rect 24574 166170 24642 166226
rect 24698 166170 24768 166226
rect 24448 166102 24768 166170
rect 24448 166046 24518 166102
rect 24574 166046 24642 166102
rect 24698 166046 24768 166102
rect 24448 165978 24768 166046
rect 24448 165922 24518 165978
rect 24574 165922 24642 165978
rect 24698 165922 24768 165978
rect 24448 165888 24768 165922
rect 55168 166350 55488 166384
rect 55168 166294 55238 166350
rect 55294 166294 55362 166350
rect 55418 166294 55488 166350
rect 55168 166226 55488 166294
rect 55168 166170 55238 166226
rect 55294 166170 55362 166226
rect 55418 166170 55488 166226
rect 55168 166102 55488 166170
rect 55168 166046 55238 166102
rect 55294 166046 55362 166102
rect 55418 166046 55488 166102
rect 55168 165978 55488 166046
rect 55168 165922 55238 165978
rect 55294 165922 55362 165978
rect 55418 165922 55488 165978
rect 55168 165888 55488 165922
rect 85888 166350 86208 166384
rect 85888 166294 85958 166350
rect 86014 166294 86082 166350
rect 86138 166294 86208 166350
rect 85888 166226 86208 166294
rect 85888 166170 85958 166226
rect 86014 166170 86082 166226
rect 86138 166170 86208 166226
rect 85888 166102 86208 166170
rect 85888 166046 85958 166102
rect 86014 166046 86082 166102
rect 86138 166046 86208 166102
rect 85888 165978 86208 166046
rect 85888 165922 85958 165978
rect 86014 165922 86082 165978
rect 86138 165922 86208 165978
rect 85888 165888 86208 165922
rect 116608 166350 116928 166384
rect 116608 166294 116678 166350
rect 116734 166294 116802 166350
rect 116858 166294 116928 166350
rect 116608 166226 116928 166294
rect 116608 166170 116678 166226
rect 116734 166170 116802 166226
rect 116858 166170 116928 166226
rect 116608 166102 116928 166170
rect 116608 166046 116678 166102
rect 116734 166046 116802 166102
rect 116858 166046 116928 166102
rect 116608 165978 116928 166046
rect 116608 165922 116678 165978
rect 116734 165922 116802 165978
rect 116858 165922 116928 165978
rect 116608 165888 116928 165922
rect 147328 166350 147648 166384
rect 147328 166294 147398 166350
rect 147454 166294 147522 166350
rect 147578 166294 147648 166350
rect 147328 166226 147648 166294
rect 147328 166170 147398 166226
rect 147454 166170 147522 166226
rect 147578 166170 147648 166226
rect 147328 166102 147648 166170
rect 147328 166046 147398 166102
rect 147454 166046 147522 166102
rect 147578 166046 147648 166102
rect 147328 165978 147648 166046
rect 147328 165922 147398 165978
rect 147454 165922 147522 165978
rect 147578 165922 147648 165978
rect 147328 165888 147648 165922
rect 178048 166350 178368 166384
rect 178048 166294 178118 166350
rect 178174 166294 178242 166350
rect 178298 166294 178368 166350
rect 178048 166226 178368 166294
rect 178048 166170 178118 166226
rect 178174 166170 178242 166226
rect 178298 166170 178368 166226
rect 178048 166102 178368 166170
rect 178048 166046 178118 166102
rect 178174 166046 178242 166102
rect 178298 166046 178368 166102
rect 178048 165978 178368 166046
rect 178048 165922 178118 165978
rect 178174 165922 178242 165978
rect 178298 165922 178368 165978
rect 178048 165888 178368 165922
rect 208768 166350 209088 166384
rect 208768 166294 208838 166350
rect 208894 166294 208962 166350
rect 209018 166294 209088 166350
rect 208768 166226 209088 166294
rect 208768 166170 208838 166226
rect 208894 166170 208962 166226
rect 209018 166170 209088 166226
rect 208768 166102 209088 166170
rect 208768 166046 208838 166102
rect 208894 166046 208962 166102
rect 209018 166046 209088 166102
rect 208768 165978 209088 166046
rect 208768 165922 208838 165978
rect 208894 165922 208962 165978
rect 209018 165922 209088 165978
rect 208768 165888 209088 165922
rect 239488 166350 239808 166384
rect 239488 166294 239558 166350
rect 239614 166294 239682 166350
rect 239738 166294 239808 166350
rect 239488 166226 239808 166294
rect 239488 166170 239558 166226
rect 239614 166170 239682 166226
rect 239738 166170 239808 166226
rect 239488 166102 239808 166170
rect 239488 166046 239558 166102
rect 239614 166046 239682 166102
rect 239738 166046 239808 166102
rect 239488 165978 239808 166046
rect 239488 165922 239558 165978
rect 239614 165922 239682 165978
rect 239738 165922 239808 165978
rect 239488 165888 239808 165922
rect 270208 166350 270528 166384
rect 270208 166294 270278 166350
rect 270334 166294 270402 166350
rect 270458 166294 270528 166350
rect 270208 166226 270528 166294
rect 270208 166170 270278 166226
rect 270334 166170 270402 166226
rect 270458 166170 270528 166226
rect 270208 166102 270528 166170
rect 270208 166046 270278 166102
rect 270334 166046 270402 166102
rect 270458 166046 270528 166102
rect 270208 165978 270528 166046
rect 270208 165922 270278 165978
rect 270334 165922 270402 165978
rect 270458 165922 270528 165978
rect 270208 165888 270528 165922
rect 300928 166350 301248 166384
rect 300928 166294 300998 166350
rect 301054 166294 301122 166350
rect 301178 166294 301248 166350
rect 300928 166226 301248 166294
rect 300928 166170 300998 166226
rect 301054 166170 301122 166226
rect 301178 166170 301248 166226
rect 300928 166102 301248 166170
rect 300928 166046 300998 166102
rect 301054 166046 301122 166102
rect 301178 166046 301248 166102
rect 300928 165978 301248 166046
rect 300928 165922 300998 165978
rect 301054 165922 301122 165978
rect 301178 165922 301248 165978
rect 300928 165888 301248 165922
rect 331648 166350 331968 166384
rect 331648 166294 331718 166350
rect 331774 166294 331842 166350
rect 331898 166294 331968 166350
rect 331648 166226 331968 166294
rect 331648 166170 331718 166226
rect 331774 166170 331842 166226
rect 331898 166170 331968 166226
rect 331648 166102 331968 166170
rect 331648 166046 331718 166102
rect 331774 166046 331842 166102
rect 331898 166046 331968 166102
rect 331648 165978 331968 166046
rect 331648 165922 331718 165978
rect 331774 165922 331842 165978
rect 331898 165922 331968 165978
rect 331648 165888 331968 165922
rect 362368 166350 362688 166384
rect 362368 166294 362438 166350
rect 362494 166294 362562 166350
rect 362618 166294 362688 166350
rect 362368 166226 362688 166294
rect 362368 166170 362438 166226
rect 362494 166170 362562 166226
rect 362618 166170 362688 166226
rect 362368 166102 362688 166170
rect 362368 166046 362438 166102
rect 362494 166046 362562 166102
rect 362618 166046 362688 166102
rect 362368 165978 362688 166046
rect 362368 165922 362438 165978
rect 362494 165922 362562 165978
rect 362618 165922 362688 165978
rect 362368 165888 362688 165922
rect 393088 166350 393408 166384
rect 393088 166294 393158 166350
rect 393214 166294 393282 166350
rect 393338 166294 393408 166350
rect 393088 166226 393408 166294
rect 393088 166170 393158 166226
rect 393214 166170 393282 166226
rect 393338 166170 393408 166226
rect 393088 166102 393408 166170
rect 393088 166046 393158 166102
rect 393214 166046 393282 166102
rect 393338 166046 393408 166102
rect 393088 165978 393408 166046
rect 393088 165922 393158 165978
rect 393214 165922 393282 165978
rect 393338 165922 393408 165978
rect 393088 165888 393408 165922
rect 423808 166350 424128 166384
rect 423808 166294 423878 166350
rect 423934 166294 424002 166350
rect 424058 166294 424128 166350
rect 423808 166226 424128 166294
rect 423808 166170 423878 166226
rect 423934 166170 424002 166226
rect 424058 166170 424128 166226
rect 423808 166102 424128 166170
rect 423808 166046 423878 166102
rect 423934 166046 424002 166102
rect 424058 166046 424128 166102
rect 423808 165978 424128 166046
rect 423808 165922 423878 165978
rect 423934 165922 424002 165978
rect 424058 165922 424128 165978
rect 423808 165888 424128 165922
rect 454528 166350 454848 166384
rect 454528 166294 454598 166350
rect 454654 166294 454722 166350
rect 454778 166294 454848 166350
rect 454528 166226 454848 166294
rect 454528 166170 454598 166226
rect 454654 166170 454722 166226
rect 454778 166170 454848 166226
rect 454528 166102 454848 166170
rect 454528 166046 454598 166102
rect 454654 166046 454722 166102
rect 454778 166046 454848 166102
rect 454528 165978 454848 166046
rect 454528 165922 454598 165978
rect 454654 165922 454722 165978
rect 454778 165922 454848 165978
rect 454528 165888 454848 165922
rect 485248 166350 485568 166384
rect 485248 166294 485318 166350
rect 485374 166294 485442 166350
rect 485498 166294 485568 166350
rect 485248 166226 485568 166294
rect 485248 166170 485318 166226
rect 485374 166170 485442 166226
rect 485498 166170 485568 166226
rect 485248 166102 485568 166170
rect 485248 166046 485318 166102
rect 485374 166046 485442 166102
rect 485498 166046 485568 166102
rect 485248 165978 485568 166046
rect 485248 165922 485318 165978
rect 485374 165922 485442 165978
rect 485498 165922 485568 165978
rect 485248 165888 485568 165922
rect 515968 166350 516288 166384
rect 515968 166294 516038 166350
rect 516094 166294 516162 166350
rect 516218 166294 516288 166350
rect 515968 166226 516288 166294
rect 515968 166170 516038 166226
rect 516094 166170 516162 166226
rect 516218 166170 516288 166226
rect 515968 166102 516288 166170
rect 515968 166046 516038 166102
rect 516094 166046 516162 166102
rect 516218 166046 516288 166102
rect 515968 165978 516288 166046
rect 515968 165922 516038 165978
rect 516094 165922 516162 165978
rect 516218 165922 516288 165978
rect 515968 165888 516288 165922
rect 525154 166350 525774 183922
rect 525154 166294 525250 166350
rect 525306 166294 525374 166350
rect 525430 166294 525498 166350
rect 525554 166294 525622 166350
rect 525678 166294 525774 166350
rect 525154 166226 525774 166294
rect 525154 166170 525250 166226
rect 525306 166170 525374 166226
rect 525430 166170 525498 166226
rect 525554 166170 525622 166226
rect 525678 166170 525774 166226
rect 525154 166102 525774 166170
rect 525154 166046 525250 166102
rect 525306 166046 525374 166102
rect 525430 166046 525498 166102
rect 525554 166046 525622 166102
rect 525678 166046 525774 166102
rect 525154 165978 525774 166046
rect 525154 165922 525250 165978
rect 525306 165922 525374 165978
rect 525430 165922 525498 165978
rect 525554 165922 525622 165978
rect 525678 165922 525774 165978
rect 6874 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 7494 154350
rect 6874 154226 7494 154294
rect 6874 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 7494 154226
rect 6874 154102 7494 154170
rect 6874 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 7494 154102
rect 6874 153978 7494 154046
rect 6874 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 7494 153978
rect 6874 136350 7494 153922
rect 39808 154350 40128 154384
rect 39808 154294 39878 154350
rect 39934 154294 40002 154350
rect 40058 154294 40128 154350
rect 39808 154226 40128 154294
rect 39808 154170 39878 154226
rect 39934 154170 40002 154226
rect 40058 154170 40128 154226
rect 39808 154102 40128 154170
rect 39808 154046 39878 154102
rect 39934 154046 40002 154102
rect 40058 154046 40128 154102
rect 39808 153978 40128 154046
rect 39808 153922 39878 153978
rect 39934 153922 40002 153978
rect 40058 153922 40128 153978
rect 39808 153888 40128 153922
rect 70528 154350 70848 154384
rect 70528 154294 70598 154350
rect 70654 154294 70722 154350
rect 70778 154294 70848 154350
rect 70528 154226 70848 154294
rect 70528 154170 70598 154226
rect 70654 154170 70722 154226
rect 70778 154170 70848 154226
rect 70528 154102 70848 154170
rect 70528 154046 70598 154102
rect 70654 154046 70722 154102
rect 70778 154046 70848 154102
rect 70528 153978 70848 154046
rect 70528 153922 70598 153978
rect 70654 153922 70722 153978
rect 70778 153922 70848 153978
rect 70528 153888 70848 153922
rect 101248 154350 101568 154384
rect 101248 154294 101318 154350
rect 101374 154294 101442 154350
rect 101498 154294 101568 154350
rect 101248 154226 101568 154294
rect 101248 154170 101318 154226
rect 101374 154170 101442 154226
rect 101498 154170 101568 154226
rect 101248 154102 101568 154170
rect 101248 154046 101318 154102
rect 101374 154046 101442 154102
rect 101498 154046 101568 154102
rect 101248 153978 101568 154046
rect 101248 153922 101318 153978
rect 101374 153922 101442 153978
rect 101498 153922 101568 153978
rect 101248 153888 101568 153922
rect 131968 154350 132288 154384
rect 131968 154294 132038 154350
rect 132094 154294 132162 154350
rect 132218 154294 132288 154350
rect 131968 154226 132288 154294
rect 131968 154170 132038 154226
rect 132094 154170 132162 154226
rect 132218 154170 132288 154226
rect 131968 154102 132288 154170
rect 131968 154046 132038 154102
rect 132094 154046 132162 154102
rect 132218 154046 132288 154102
rect 131968 153978 132288 154046
rect 131968 153922 132038 153978
rect 132094 153922 132162 153978
rect 132218 153922 132288 153978
rect 131968 153888 132288 153922
rect 162688 154350 163008 154384
rect 162688 154294 162758 154350
rect 162814 154294 162882 154350
rect 162938 154294 163008 154350
rect 162688 154226 163008 154294
rect 162688 154170 162758 154226
rect 162814 154170 162882 154226
rect 162938 154170 163008 154226
rect 162688 154102 163008 154170
rect 162688 154046 162758 154102
rect 162814 154046 162882 154102
rect 162938 154046 163008 154102
rect 162688 153978 163008 154046
rect 162688 153922 162758 153978
rect 162814 153922 162882 153978
rect 162938 153922 163008 153978
rect 162688 153888 163008 153922
rect 193408 154350 193728 154384
rect 193408 154294 193478 154350
rect 193534 154294 193602 154350
rect 193658 154294 193728 154350
rect 193408 154226 193728 154294
rect 193408 154170 193478 154226
rect 193534 154170 193602 154226
rect 193658 154170 193728 154226
rect 193408 154102 193728 154170
rect 193408 154046 193478 154102
rect 193534 154046 193602 154102
rect 193658 154046 193728 154102
rect 193408 153978 193728 154046
rect 193408 153922 193478 153978
rect 193534 153922 193602 153978
rect 193658 153922 193728 153978
rect 193408 153888 193728 153922
rect 224128 154350 224448 154384
rect 224128 154294 224198 154350
rect 224254 154294 224322 154350
rect 224378 154294 224448 154350
rect 224128 154226 224448 154294
rect 224128 154170 224198 154226
rect 224254 154170 224322 154226
rect 224378 154170 224448 154226
rect 224128 154102 224448 154170
rect 224128 154046 224198 154102
rect 224254 154046 224322 154102
rect 224378 154046 224448 154102
rect 224128 153978 224448 154046
rect 224128 153922 224198 153978
rect 224254 153922 224322 153978
rect 224378 153922 224448 153978
rect 224128 153888 224448 153922
rect 254848 154350 255168 154384
rect 254848 154294 254918 154350
rect 254974 154294 255042 154350
rect 255098 154294 255168 154350
rect 254848 154226 255168 154294
rect 254848 154170 254918 154226
rect 254974 154170 255042 154226
rect 255098 154170 255168 154226
rect 254848 154102 255168 154170
rect 254848 154046 254918 154102
rect 254974 154046 255042 154102
rect 255098 154046 255168 154102
rect 254848 153978 255168 154046
rect 254848 153922 254918 153978
rect 254974 153922 255042 153978
rect 255098 153922 255168 153978
rect 254848 153888 255168 153922
rect 285568 154350 285888 154384
rect 285568 154294 285638 154350
rect 285694 154294 285762 154350
rect 285818 154294 285888 154350
rect 285568 154226 285888 154294
rect 285568 154170 285638 154226
rect 285694 154170 285762 154226
rect 285818 154170 285888 154226
rect 285568 154102 285888 154170
rect 285568 154046 285638 154102
rect 285694 154046 285762 154102
rect 285818 154046 285888 154102
rect 285568 153978 285888 154046
rect 285568 153922 285638 153978
rect 285694 153922 285762 153978
rect 285818 153922 285888 153978
rect 285568 153888 285888 153922
rect 316288 154350 316608 154384
rect 316288 154294 316358 154350
rect 316414 154294 316482 154350
rect 316538 154294 316608 154350
rect 316288 154226 316608 154294
rect 316288 154170 316358 154226
rect 316414 154170 316482 154226
rect 316538 154170 316608 154226
rect 316288 154102 316608 154170
rect 316288 154046 316358 154102
rect 316414 154046 316482 154102
rect 316538 154046 316608 154102
rect 316288 153978 316608 154046
rect 316288 153922 316358 153978
rect 316414 153922 316482 153978
rect 316538 153922 316608 153978
rect 316288 153888 316608 153922
rect 347008 154350 347328 154384
rect 347008 154294 347078 154350
rect 347134 154294 347202 154350
rect 347258 154294 347328 154350
rect 347008 154226 347328 154294
rect 347008 154170 347078 154226
rect 347134 154170 347202 154226
rect 347258 154170 347328 154226
rect 347008 154102 347328 154170
rect 347008 154046 347078 154102
rect 347134 154046 347202 154102
rect 347258 154046 347328 154102
rect 347008 153978 347328 154046
rect 347008 153922 347078 153978
rect 347134 153922 347202 153978
rect 347258 153922 347328 153978
rect 347008 153888 347328 153922
rect 377728 154350 378048 154384
rect 377728 154294 377798 154350
rect 377854 154294 377922 154350
rect 377978 154294 378048 154350
rect 377728 154226 378048 154294
rect 377728 154170 377798 154226
rect 377854 154170 377922 154226
rect 377978 154170 378048 154226
rect 377728 154102 378048 154170
rect 377728 154046 377798 154102
rect 377854 154046 377922 154102
rect 377978 154046 378048 154102
rect 377728 153978 378048 154046
rect 377728 153922 377798 153978
rect 377854 153922 377922 153978
rect 377978 153922 378048 153978
rect 377728 153888 378048 153922
rect 408448 154350 408768 154384
rect 408448 154294 408518 154350
rect 408574 154294 408642 154350
rect 408698 154294 408768 154350
rect 408448 154226 408768 154294
rect 408448 154170 408518 154226
rect 408574 154170 408642 154226
rect 408698 154170 408768 154226
rect 408448 154102 408768 154170
rect 408448 154046 408518 154102
rect 408574 154046 408642 154102
rect 408698 154046 408768 154102
rect 408448 153978 408768 154046
rect 408448 153922 408518 153978
rect 408574 153922 408642 153978
rect 408698 153922 408768 153978
rect 408448 153888 408768 153922
rect 439168 154350 439488 154384
rect 439168 154294 439238 154350
rect 439294 154294 439362 154350
rect 439418 154294 439488 154350
rect 439168 154226 439488 154294
rect 439168 154170 439238 154226
rect 439294 154170 439362 154226
rect 439418 154170 439488 154226
rect 439168 154102 439488 154170
rect 439168 154046 439238 154102
rect 439294 154046 439362 154102
rect 439418 154046 439488 154102
rect 439168 153978 439488 154046
rect 439168 153922 439238 153978
rect 439294 153922 439362 153978
rect 439418 153922 439488 153978
rect 439168 153888 439488 153922
rect 469888 154350 470208 154384
rect 469888 154294 469958 154350
rect 470014 154294 470082 154350
rect 470138 154294 470208 154350
rect 469888 154226 470208 154294
rect 469888 154170 469958 154226
rect 470014 154170 470082 154226
rect 470138 154170 470208 154226
rect 469888 154102 470208 154170
rect 469888 154046 469958 154102
rect 470014 154046 470082 154102
rect 470138 154046 470208 154102
rect 469888 153978 470208 154046
rect 469888 153922 469958 153978
rect 470014 153922 470082 153978
rect 470138 153922 470208 153978
rect 469888 153888 470208 153922
rect 500608 154350 500928 154384
rect 500608 154294 500678 154350
rect 500734 154294 500802 154350
rect 500858 154294 500928 154350
rect 500608 154226 500928 154294
rect 500608 154170 500678 154226
rect 500734 154170 500802 154226
rect 500858 154170 500928 154226
rect 500608 154102 500928 154170
rect 500608 154046 500678 154102
rect 500734 154046 500802 154102
rect 500858 154046 500928 154102
rect 500608 153978 500928 154046
rect 500608 153922 500678 153978
rect 500734 153922 500802 153978
rect 500858 153922 500928 153978
rect 500608 153888 500928 153922
rect 24448 148350 24768 148384
rect 24448 148294 24518 148350
rect 24574 148294 24642 148350
rect 24698 148294 24768 148350
rect 24448 148226 24768 148294
rect 24448 148170 24518 148226
rect 24574 148170 24642 148226
rect 24698 148170 24768 148226
rect 24448 148102 24768 148170
rect 24448 148046 24518 148102
rect 24574 148046 24642 148102
rect 24698 148046 24768 148102
rect 24448 147978 24768 148046
rect 24448 147922 24518 147978
rect 24574 147922 24642 147978
rect 24698 147922 24768 147978
rect 24448 147888 24768 147922
rect 55168 148350 55488 148384
rect 55168 148294 55238 148350
rect 55294 148294 55362 148350
rect 55418 148294 55488 148350
rect 55168 148226 55488 148294
rect 55168 148170 55238 148226
rect 55294 148170 55362 148226
rect 55418 148170 55488 148226
rect 55168 148102 55488 148170
rect 55168 148046 55238 148102
rect 55294 148046 55362 148102
rect 55418 148046 55488 148102
rect 55168 147978 55488 148046
rect 55168 147922 55238 147978
rect 55294 147922 55362 147978
rect 55418 147922 55488 147978
rect 55168 147888 55488 147922
rect 85888 148350 86208 148384
rect 85888 148294 85958 148350
rect 86014 148294 86082 148350
rect 86138 148294 86208 148350
rect 85888 148226 86208 148294
rect 85888 148170 85958 148226
rect 86014 148170 86082 148226
rect 86138 148170 86208 148226
rect 85888 148102 86208 148170
rect 85888 148046 85958 148102
rect 86014 148046 86082 148102
rect 86138 148046 86208 148102
rect 85888 147978 86208 148046
rect 85888 147922 85958 147978
rect 86014 147922 86082 147978
rect 86138 147922 86208 147978
rect 85888 147888 86208 147922
rect 116608 148350 116928 148384
rect 116608 148294 116678 148350
rect 116734 148294 116802 148350
rect 116858 148294 116928 148350
rect 116608 148226 116928 148294
rect 116608 148170 116678 148226
rect 116734 148170 116802 148226
rect 116858 148170 116928 148226
rect 116608 148102 116928 148170
rect 116608 148046 116678 148102
rect 116734 148046 116802 148102
rect 116858 148046 116928 148102
rect 116608 147978 116928 148046
rect 116608 147922 116678 147978
rect 116734 147922 116802 147978
rect 116858 147922 116928 147978
rect 116608 147888 116928 147922
rect 147328 148350 147648 148384
rect 147328 148294 147398 148350
rect 147454 148294 147522 148350
rect 147578 148294 147648 148350
rect 147328 148226 147648 148294
rect 147328 148170 147398 148226
rect 147454 148170 147522 148226
rect 147578 148170 147648 148226
rect 147328 148102 147648 148170
rect 147328 148046 147398 148102
rect 147454 148046 147522 148102
rect 147578 148046 147648 148102
rect 147328 147978 147648 148046
rect 147328 147922 147398 147978
rect 147454 147922 147522 147978
rect 147578 147922 147648 147978
rect 147328 147888 147648 147922
rect 178048 148350 178368 148384
rect 178048 148294 178118 148350
rect 178174 148294 178242 148350
rect 178298 148294 178368 148350
rect 178048 148226 178368 148294
rect 178048 148170 178118 148226
rect 178174 148170 178242 148226
rect 178298 148170 178368 148226
rect 178048 148102 178368 148170
rect 178048 148046 178118 148102
rect 178174 148046 178242 148102
rect 178298 148046 178368 148102
rect 178048 147978 178368 148046
rect 178048 147922 178118 147978
rect 178174 147922 178242 147978
rect 178298 147922 178368 147978
rect 178048 147888 178368 147922
rect 208768 148350 209088 148384
rect 208768 148294 208838 148350
rect 208894 148294 208962 148350
rect 209018 148294 209088 148350
rect 208768 148226 209088 148294
rect 208768 148170 208838 148226
rect 208894 148170 208962 148226
rect 209018 148170 209088 148226
rect 208768 148102 209088 148170
rect 208768 148046 208838 148102
rect 208894 148046 208962 148102
rect 209018 148046 209088 148102
rect 208768 147978 209088 148046
rect 208768 147922 208838 147978
rect 208894 147922 208962 147978
rect 209018 147922 209088 147978
rect 208768 147888 209088 147922
rect 239488 148350 239808 148384
rect 239488 148294 239558 148350
rect 239614 148294 239682 148350
rect 239738 148294 239808 148350
rect 239488 148226 239808 148294
rect 239488 148170 239558 148226
rect 239614 148170 239682 148226
rect 239738 148170 239808 148226
rect 239488 148102 239808 148170
rect 239488 148046 239558 148102
rect 239614 148046 239682 148102
rect 239738 148046 239808 148102
rect 239488 147978 239808 148046
rect 239488 147922 239558 147978
rect 239614 147922 239682 147978
rect 239738 147922 239808 147978
rect 239488 147888 239808 147922
rect 270208 148350 270528 148384
rect 270208 148294 270278 148350
rect 270334 148294 270402 148350
rect 270458 148294 270528 148350
rect 270208 148226 270528 148294
rect 270208 148170 270278 148226
rect 270334 148170 270402 148226
rect 270458 148170 270528 148226
rect 270208 148102 270528 148170
rect 270208 148046 270278 148102
rect 270334 148046 270402 148102
rect 270458 148046 270528 148102
rect 270208 147978 270528 148046
rect 270208 147922 270278 147978
rect 270334 147922 270402 147978
rect 270458 147922 270528 147978
rect 270208 147888 270528 147922
rect 300928 148350 301248 148384
rect 300928 148294 300998 148350
rect 301054 148294 301122 148350
rect 301178 148294 301248 148350
rect 300928 148226 301248 148294
rect 300928 148170 300998 148226
rect 301054 148170 301122 148226
rect 301178 148170 301248 148226
rect 300928 148102 301248 148170
rect 300928 148046 300998 148102
rect 301054 148046 301122 148102
rect 301178 148046 301248 148102
rect 300928 147978 301248 148046
rect 300928 147922 300998 147978
rect 301054 147922 301122 147978
rect 301178 147922 301248 147978
rect 300928 147888 301248 147922
rect 331648 148350 331968 148384
rect 331648 148294 331718 148350
rect 331774 148294 331842 148350
rect 331898 148294 331968 148350
rect 331648 148226 331968 148294
rect 331648 148170 331718 148226
rect 331774 148170 331842 148226
rect 331898 148170 331968 148226
rect 331648 148102 331968 148170
rect 331648 148046 331718 148102
rect 331774 148046 331842 148102
rect 331898 148046 331968 148102
rect 331648 147978 331968 148046
rect 331648 147922 331718 147978
rect 331774 147922 331842 147978
rect 331898 147922 331968 147978
rect 331648 147888 331968 147922
rect 362368 148350 362688 148384
rect 362368 148294 362438 148350
rect 362494 148294 362562 148350
rect 362618 148294 362688 148350
rect 362368 148226 362688 148294
rect 362368 148170 362438 148226
rect 362494 148170 362562 148226
rect 362618 148170 362688 148226
rect 362368 148102 362688 148170
rect 362368 148046 362438 148102
rect 362494 148046 362562 148102
rect 362618 148046 362688 148102
rect 362368 147978 362688 148046
rect 362368 147922 362438 147978
rect 362494 147922 362562 147978
rect 362618 147922 362688 147978
rect 362368 147888 362688 147922
rect 393088 148350 393408 148384
rect 393088 148294 393158 148350
rect 393214 148294 393282 148350
rect 393338 148294 393408 148350
rect 393088 148226 393408 148294
rect 393088 148170 393158 148226
rect 393214 148170 393282 148226
rect 393338 148170 393408 148226
rect 393088 148102 393408 148170
rect 393088 148046 393158 148102
rect 393214 148046 393282 148102
rect 393338 148046 393408 148102
rect 393088 147978 393408 148046
rect 393088 147922 393158 147978
rect 393214 147922 393282 147978
rect 393338 147922 393408 147978
rect 393088 147888 393408 147922
rect 423808 148350 424128 148384
rect 423808 148294 423878 148350
rect 423934 148294 424002 148350
rect 424058 148294 424128 148350
rect 423808 148226 424128 148294
rect 423808 148170 423878 148226
rect 423934 148170 424002 148226
rect 424058 148170 424128 148226
rect 423808 148102 424128 148170
rect 423808 148046 423878 148102
rect 423934 148046 424002 148102
rect 424058 148046 424128 148102
rect 423808 147978 424128 148046
rect 423808 147922 423878 147978
rect 423934 147922 424002 147978
rect 424058 147922 424128 147978
rect 423808 147888 424128 147922
rect 454528 148350 454848 148384
rect 454528 148294 454598 148350
rect 454654 148294 454722 148350
rect 454778 148294 454848 148350
rect 454528 148226 454848 148294
rect 454528 148170 454598 148226
rect 454654 148170 454722 148226
rect 454778 148170 454848 148226
rect 454528 148102 454848 148170
rect 454528 148046 454598 148102
rect 454654 148046 454722 148102
rect 454778 148046 454848 148102
rect 454528 147978 454848 148046
rect 454528 147922 454598 147978
rect 454654 147922 454722 147978
rect 454778 147922 454848 147978
rect 454528 147888 454848 147922
rect 485248 148350 485568 148384
rect 485248 148294 485318 148350
rect 485374 148294 485442 148350
rect 485498 148294 485568 148350
rect 485248 148226 485568 148294
rect 485248 148170 485318 148226
rect 485374 148170 485442 148226
rect 485498 148170 485568 148226
rect 485248 148102 485568 148170
rect 485248 148046 485318 148102
rect 485374 148046 485442 148102
rect 485498 148046 485568 148102
rect 485248 147978 485568 148046
rect 485248 147922 485318 147978
rect 485374 147922 485442 147978
rect 485498 147922 485568 147978
rect 485248 147888 485568 147922
rect 515968 148350 516288 148384
rect 515968 148294 516038 148350
rect 516094 148294 516162 148350
rect 516218 148294 516288 148350
rect 515968 148226 516288 148294
rect 515968 148170 516038 148226
rect 516094 148170 516162 148226
rect 516218 148170 516288 148226
rect 515968 148102 516288 148170
rect 515968 148046 516038 148102
rect 516094 148046 516162 148102
rect 516218 148046 516288 148102
rect 515968 147978 516288 148046
rect 515968 147922 516038 147978
rect 516094 147922 516162 147978
rect 516218 147922 516288 147978
rect 515968 147888 516288 147922
rect 525154 148350 525774 165922
rect 525154 148294 525250 148350
rect 525306 148294 525374 148350
rect 525430 148294 525498 148350
rect 525554 148294 525622 148350
rect 525678 148294 525774 148350
rect 525154 148226 525774 148294
rect 525154 148170 525250 148226
rect 525306 148170 525374 148226
rect 525430 148170 525498 148226
rect 525554 148170 525622 148226
rect 525678 148170 525774 148226
rect 525154 148102 525774 148170
rect 525154 148046 525250 148102
rect 525306 148046 525374 148102
rect 525430 148046 525498 148102
rect 525554 148046 525622 148102
rect 525678 148046 525774 148102
rect 525154 147978 525774 148046
rect 525154 147922 525250 147978
rect 525306 147922 525374 147978
rect 525430 147922 525498 147978
rect 525554 147922 525622 147978
rect 525678 147922 525774 147978
rect 6874 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 7494 136350
rect 6874 136226 7494 136294
rect 6874 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 7494 136226
rect 6874 136102 7494 136170
rect 6874 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 7494 136102
rect 6874 135978 7494 136046
rect 6874 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 7494 135978
rect 6874 118350 7494 135922
rect 39808 136350 40128 136384
rect 39808 136294 39878 136350
rect 39934 136294 40002 136350
rect 40058 136294 40128 136350
rect 39808 136226 40128 136294
rect 39808 136170 39878 136226
rect 39934 136170 40002 136226
rect 40058 136170 40128 136226
rect 39808 136102 40128 136170
rect 39808 136046 39878 136102
rect 39934 136046 40002 136102
rect 40058 136046 40128 136102
rect 39808 135978 40128 136046
rect 39808 135922 39878 135978
rect 39934 135922 40002 135978
rect 40058 135922 40128 135978
rect 39808 135888 40128 135922
rect 70528 136350 70848 136384
rect 70528 136294 70598 136350
rect 70654 136294 70722 136350
rect 70778 136294 70848 136350
rect 70528 136226 70848 136294
rect 70528 136170 70598 136226
rect 70654 136170 70722 136226
rect 70778 136170 70848 136226
rect 70528 136102 70848 136170
rect 70528 136046 70598 136102
rect 70654 136046 70722 136102
rect 70778 136046 70848 136102
rect 70528 135978 70848 136046
rect 70528 135922 70598 135978
rect 70654 135922 70722 135978
rect 70778 135922 70848 135978
rect 70528 135888 70848 135922
rect 101248 136350 101568 136384
rect 101248 136294 101318 136350
rect 101374 136294 101442 136350
rect 101498 136294 101568 136350
rect 101248 136226 101568 136294
rect 101248 136170 101318 136226
rect 101374 136170 101442 136226
rect 101498 136170 101568 136226
rect 101248 136102 101568 136170
rect 101248 136046 101318 136102
rect 101374 136046 101442 136102
rect 101498 136046 101568 136102
rect 101248 135978 101568 136046
rect 101248 135922 101318 135978
rect 101374 135922 101442 135978
rect 101498 135922 101568 135978
rect 101248 135888 101568 135922
rect 131968 136350 132288 136384
rect 131968 136294 132038 136350
rect 132094 136294 132162 136350
rect 132218 136294 132288 136350
rect 131968 136226 132288 136294
rect 131968 136170 132038 136226
rect 132094 136170 132162 136226
rect 132218 136170 132288 136226
rect 131968 136102 132288 136170
rect 131968 136046 132038 136102
rect 132094 136046 132162 136102
rect 132218 136046 132288 136102
rect 131968 135978 132288 136046
rect 131968 135922 132038 135978
rect 132094 135922 132162 135978
rect 132218 135922 132288 135978
rect 131968 135888 132288 135922
rect 162688 136350 163008 136384
rect 162688 136294 162758 136350
rect 162814 136294 162882 136350
rect 162938 136294 163008 136350
rect 162688 136226 163008 136294
rect 162688 136170 162758 136226
rect 162814 136170 162882 136226
rect 162938 136170 163008 136226
rect 162688 136102 163008 136170
rect 162688 136046 162758 136102
rect 162814 136046 162882 136102
rect 162938 136046 163008 136102
rect 162688 135978 163008 136046
rect 162688 135922 162758 135978
rect 162814 135922 162882 135978
rect 162938 135922 163008 135978
rect 162688 135888 163008 135922
rect 193408 136350 193728 136384
rect 193408 136294 193478 136350
rect 193534 136294 193602 136350
rect 193658 136294 193728 136350
rect 193408 136226 193728 136294
rect 193408 136170 193478 136226
rect 193534 136170 193602 136226
rect 193658 136170 193728 136226
rect 193408 136102 193728 136170
rect 193408 136046 193478 136102
rect 193534 136046 193602 136102
rect 193658 136046 193728 136102
rect 193408 135978 193728 136046
rect 193408 135922 193478 135978
rect 193534 135922 193602 135978
rect 193658 135922 193728 135978
rect 193408 135888 193728 135922
rect 224128 136350 224448 136384
rect 224128 136294 224198 136350
rect 224254 136294 224322 136350
rect 224378 136294 224448 136350
rect 224128 136226 224448 136294
rect 224128 136170 224198 136226
rect 224254 136170 224322 136226
rect 224378 136170 224448 136226
rect 224128 136102 224448 136170
rect 224128 136046 224198 136102
rect 224254 136046 224322 136102
rect 224378 136046 224448 136102
rect 224128 135978 224448 136046
rect 224128 135922 224198 135978
rect 224254 135922 224322 135978
rect 224378 135922 224448 135978
rect 224128 135888 224448 135922
rect 254848 136350 255168 136384
rect 254848 136294 254918 136350
rect 254974 136294 255042 136350
rect 255098 136294 255168 136350
rect 254848 136226 255168 136294
rect 254848 136170 254918 136226
rect 254974 136170 255042 136226
rect 255098 136170 255168 136226
rect 254848 136102 255168 136170
rect 254848 136046 254918 136102
rect 254974 136046 255042 136102
rect 255098 136046 255168 136102
rect 254848 135978 255168 136046
rect 254848 135922 254918 135978
rect 254974 135922 255042 135978
rect 255098 135922 255168 135978
rect 254848 135888 255168 135922
rect 285568 136350 285888 136384
rect 285568 136294 285638 136350
rect 285694 136294 285762 136350
rect 285818 136294 285888 136350
rect 285568 136226 285888 136294
rect 285568 136170 285638 136226
rect 285694 136170 285762 136226
rect 285818 136170 285888 136226
rect 285568 136102 285888 136170
rect 285568 136046 285638 136102
rect 285694 136046 285762 136102
rect 285818 136046 285888 136102
rect 285568 135978 285888 136046
rect 285568 135922 285638 135978
rect 285694 135922 285762 135978
rect 285818 135922 285888 135978
rect 285568 135888 285888 135922
rect 316288 136350 316608 136384
rect 316288 136294 316358 136350
rect 316414 136294 316482 136350
rect 316538 136294 316608 136350
rect 316288 136226 316608 136294
rect 316288 136170 316358 136226
rect 316414 136170 316482 136226
rect 316538 136170 316608 136226
rect 316288 136102 316608 136170
rect 316288 136046 316358 136102
rect 316414 136046 316482 136102
rect 316538 136046 316608 136102
rect 316288 135978 316608 136046
rect 316288 135922 316358 135978
rect 316414 135922 316482 135978
rect 316538 135922 316608 135978
rect 316288 135888 316608 135922
rect 347008 136350 347328 136384
rect 347008 136294 347078 136350
rect 347134 136294 347202 136350
rect 347258 136294 347328 136350
rect 347008 136226 347328 136294
rect 347008 136170 347078 136226
rect 347134 136170 347202 136226
rect 347258 136170 347328 136226
rect 347008 136102 347328 136170
rect 347008 136046 347078 136102
rect 347134 136046 347202 136102
rect 347258 136046 347328 136102
rect 347008 135978 347328 136046
rect 347008 135922 347078 135978
rect 347134 135922 347202 135978
rect 347258 135922 347328 135978
rect 347008 135888 347328 135922
rect 377728 136350 378048 136384
rect 377728 136294 377798 136350
rect 377854 136294 377922 136350
rect 377978 136294 378048 136350
rect 377728 136226 378048 136294
rect 377728 136170 377798 136226
rect 377854 136170 377922 136226
rect 377978 136170 378048 136226
rect 377728 136102 378048 136170
rect 377728 136046 377798 136102
rect 377854 136046 377922 136102
rect 377978 136046 378048 136102
rect 377728 135978 378048 136046
rect 377728 135922 377798 135978
rect 377854 135922 377922 135978
rect 377978 135922 378048 135978
rect 377728 135888 378048 135922
rect 408448 136350 408768 136384
rect 408448 136294 408518 136350
rect 408574 136294 408642 136350
rect 408698 136294 408768 136350
rect 408448 136226 408768 136294
rect 408448 136170 408518 136226
rect 408574 136170 408642 136226
rect 408698 136170 408768 136226
rect 408448 136102 408768 136170
rect 408448 136046 408518 136102
rect 408574 136046 408642 136102
rect 408698 136046 408768 136102
rect 408448 135978 408768 136046
rect 408448 135922 408518 135978
rect 408574 135922 408642 135978
rect 408698 135922 408768 135978
rect 408448 135888 408768 135922
rect 439168 136350 439488 136384
rect 439168 136294 439238 136350
rect 439294 136294 439362 136350
rect 439418 136294 439488 136350
rect 439168 136226 439488 136294
rect 439168 136170 439238 136226
rect 439294 136170 439362 136226
rect 439418 136170 439488 136226
rect 439168 136102 439488 136170
rect 439168 136046 439238 136102
rect 439294 136046 439362 136102
rect 439418 136046 439488 136102
rect 439168 135978 439488 136046
rect 439168 135922 439238 135978
rect 439294 135922 439362 135978
rect 439418 135922 439488 135978
rect 439168 135888 439488 135922
rect 469888 136350 470208 136384
rect 469888 136294 469958 136350
rect 470014 136294 470082 136350
rect 470138 136294 470208 136350
rect 469888 136226 470208 136294
rect 469888 136170 469958 136226
rect 470014 136170 470082 136226
rect 470138 136170 470208 136226
rect 469888 136102 470208 136170
rect 469888 136046 469958 136102
rect 470014 136046 470082 136102
rect 470138 136046 470208 136102
rect 469888 135978 470208 136046
rect 469888 135922 469958 135978
rect 470014 135922 470082 135978
rect 470138 135922 470208 135978
rect 469888 135888 470208 135922
rect 500608 136350 500928 136384
rect 500608 136294 500678 136350
rect 500734 136294 500802 136350
rect 500858 136294 500928 136350
rect 500608 136226 500928 136294
rect 500608 136170 500678 136226
rect 500734 136170 500802 136226
rect 500858 136170 500928 136226
rect 500608 136102 500928 136170
rect 500608 136046 500678 136102
rect 500734 136046 500802 136102
rect 500858 136046 500928 136102
rect 500608 135978 500928 136046
rect 500608 135922 500678 135978
rect 500734 135922 500802 135978
rect 500858 135922 500928 135978
rect 500608 135888 500928 135922
rect 24448 130350 24768 130384
rect 24448 130294 24518 130350
rect 24574 130294 24642 130350
rect 24698 130294 24768 130350
rect 24448 130226 24768 130294
rect 24448 130170 24518 130226
rect 24574 130170 24642 130226
rect 24698 130170 24768 130226
rect 24448 130102 24768 130170
rect 24448 130046 24518 130102
rect 24574 130046 24642 130102
rect 24698 130046 24768 130102
rect 24448 129978 24768 130046
rect 24448 129922 24518 129978
rect 24574 129922 24642 129978
rect 24698 129922 24768 129978
rect 24448 129888 24768 129922
rect 55168 130350 55488 130384
rect 55168 130294 55238 130350
rect 55294 130294 55362 130350
rect 55418 130294 55488 130350
rect 55168 130226 55488 130294
rect 55168 130170 55238 130226
rect 55294 130170 55362 130226
rect 55418 130170 55488 130226
rect 55168 130102 55488 130170
rect 55168 130046 55238 130102
rect 55294 130046 55362 130102
rect 55418 130046 55488 130102
rect 55168 129978 55488 130046
rect 55168 129922 55238 129978
rect 55294 129922 55362 129978
rect 55418 129922 55488 129978
rect 55168 129888 55488 129922
rect 85888 130350 86208 130384
rect 85888 130294 85958 130350
rect 86014 130294 86082 130350
rect 86138 130294 86208 130350
rect 85888 130226 86208 130294
rect 85888 130170 85958 130226
rect 86014 130170 86082 130226
rect 86138 130170 86208 130226
rect 85888 130102 86208 130170
rect 85888 130046 85958 130102
rect 86014 130046 86082 130102
rect 86138 130046 86208 130102
rect 85888 129978 86208 130046
rect 85888 129922 85958 129978
rect 86014 129922 86082 129978
rect 86138 129922 86208 129978
rect 85888 129888 86208 129922
rect 116608 130350 116928 130384
rect 116608 130294 116678 130350
rect 116734 130294 116802 130350
rect 116858 130294 116928 130350
rect 116608 130226 116928 130294
rect 116608 130170 116678 130226
rect 116734 130170 116802 130226
rect 116858 130170 116928 130226
rect 116608 130102 116928 130170
rect 116608 130046 116678 130102
rect 116734 130046 116802 130102
rect 116858 130046 116928 130102
rect 116608 129978 116928 130046
rect 116608 129922 116678 129978
rect 116734 129922 116802 129978
rect 116858 129922 116928 129978
rect 116608 129888 116928 129922
rect 147328 130350 147648 130384
rect 147328 130294 147398 130350
rect 147454 130294 147522 130350
rect 147578 130294 147648 130350
rect 147328 130226 147648 130294
rect 147328 130170 147398 130226
rect 147454 130170 147522 130226
rect 147578 130170 147648 130226
rect 147328 130102 147648 130170
rect 147328 130046 147398 130102
rect 147454 130046 147522 130102
rect 147578 130046 147648 130102
rect 147328 129978 147648 130046
rect 147328 129922 147398 129978
rect 147454 129922 147522 129978
rect 147578 129922 147648 129978
rect 147328 129888 147648 129922
rect 178048 130350 178368 130384
rect 178048 130294 178118 130350
rect 178174 130294 178242 130350
rect 178298 130294 178368 130350
rect 178048 130226 178368 130294
rect 178048 130170 178118 130226
rect 178174 130170 178242 130226
rect 178298 130170 178368 130226
rect 178048 130102 178368 130170
rect 178048 130046 178118 130102
rect 178174 130046 178242 130102
rect 178298 130046 178368 130102
rect 178048 129978 178368 130046
rect 178048 129922 178118 129978
rect 178174 129922 178242 129978
rect 178298 129922 178368 129978
rect 178048 129888 178368 129922
rect 208768 130350 209088 130384
rect 208768 130294 208838 130350
rect 208894 130294 208962 130350
rect 209018 130294 209088 130350
rect 208768 130226 209088 130294
rect 208768 130170 208838 130226
rect 208894 130170 208962 130226
rect 209018 130170 209088 130226
rect 208768 130102 209088 130170
rect 208768 130046 208838 130102
rect 208894 130046 208962 130102
rect 209018 130046 209088 130102
rect 208768 129978 209088 130046
rect 208768 129922 208838 129978
rect 208894 129922 208962 129978
rect 209018 129922 209088 129978
rect 208768 129888 209088 129922
rect 239488 130350 239808 130384
rect 239488 130294 239558 130350
rect 239614 130294 239682 130350
rect 239738 130294 239808 130350
rect 239488 130226 239808 130294
rect 239488 130170 239558 130226
rect 239614 130170 239682 130226
rect 239738 130170 239808 130226
rect 239488 130102 239808 130170
rect 239488 130046 239558 130102
rect 239614 130046 239682 130102
rect 239738 130046 239808 130102
rect 239488 129978 239808 130046
rect 239488 129922 239558 129978
rect 239614 129922 239682 129978
rect 239738 129922 239808 129978
rect 239488 129888 239808 129922
rect 270208 130350 270528 130384
rect 270208 130294 270278 130350
rect 270334 130294 270402 130350
rect 270458 130294 270528 130350
rect 270208 130226 270528 130294
rect 270208 130170 270278 130226
rect 270334 130170 270402 130226
rect 270458 130170 270528 130226
rect 270208 130102 270528 130170
rect 270208 130046 270278 130102
rect 270334 130046 270402 130102
rect 270458 130046 270528 130102
rect 270208 129978 270528 130046
rect 270208 129922 270278 129978
rect 270334 129922 270402 129978
rect 270458 129922 270528 129978
rect 270208 129888 270528 129922
rect 300928 130350 301248 130384
rect 300928 130294 300998 130350
rect 301054 130294 301122 130350
rect 301178 130294 301248 130350
rect 300928 130226 301248 130294
rect 300928 130170 300998 130226
rect 301054 130170 301122 130226
rect 301178 130170 301248 130226
rect 300928 130102 301248 130170
rect 300928 130046 300998 130102
rect 301054 130046 301122 130102
rect 301178 130046 301248 130102
rect 300928 129978 301248 130046
rect 300928 129922 300998 129978
rect 301054 129922 301122 129978
rect 301178 129922 301248 129978
rect 300928 129888 301248 129922
rect 331648 130350 331968 130384
rect 331648 130294 331718 130350
rect 331774 130294 331842 130350
rect 331898 130294 331968 130350
rect 331648 130226 331968 130294
rect 331648 130170 331718 130226
rect 331774 130170 331842 130226
rect 331898 130170 331968 130226
rect 331648 130102 331968 130170
rect 331648 130046 331718 130102
rect 331774 130046 331842 130102
rect 331898 130046 331968 130102
rect 331648 129978 331968 130046
rect 331648 129922 331718 129978
rect 331774 129922 331842 129978
rect 331898 129922 331968 129978
rect 331648 129888 331968 129922
rect 362368 130350 362688 130384
rect 362368 130294 362438 130350
rect 362494 130294 362562 130350
rect 362618 130294 362688 130350
rect 362368 130226 362688 130294
rect 362368 130170 362438 130226
rect 362494 130170 362562 130226
rect 362618 130170 362688 130226
rect 362368 130102 362688 130170
rect 362368 130046 362438 130102
rect 362494 130046 362562 130102
rect 362618 130046 362688 130102
rect 362368 129978 362688 130046
rect 362368 129922 362438 129978
rect 362494 129922 362562 129978
rect 362618 129922 362688 129978
rect 362368 129888 362688 129922
rect 393088 130350 393408 130384
rect 393088 130294 393158 130350
rect 393214 130294 393282 130350
rect 393338 130294 393408 130350
rect 393088 130226 393408 130294
rect 393088 130170 393158 130226
rect 393214 130170 393282 130226
rect 393338 130170 393408 130226
rect 393088 130102 393408 130170
rect 393088 130046 393158 130102
rect 393214 130046 393282 130102
rect 393338 130046 393408 130102
rect 393088 129978 393408 130046
rect 393088 129922 393158 129978
rect 393214 129922 393282 129978
rect 393338 129922 393408 129978
rect 393088 129888 393408 129922
rect 423808 130350 424128 130384
rect 423808 130294 423878 130350
rect 423934 130294 424002 130350
rect 424058 130294 424128 130350
rect 423808 130226 424128 130294
rect 423808 130170 423878 130226
rect 423934 130170 424002 130226
rect 424058 130170 424128 130226
rect 423808 130102 424128 130170
rect 423808 130046 423878 130102
rect 423934 130046 424002 130102
rect 424058 130046 424128 130102
rect 423808 129978 424128 130046
rect 423808 129922 423878 129978
rect 423934 129922 424002 129978
rect 424058 129922 424128 129978
rect 423808 129888 424128 129922
rect 454528 130350 454848 130384
rect 454528 130294 454598 130350
rect 454654 130294 454722 130350
rect 454778 130294 454848 130350
rect 454528 130226 454848 130294
rect 454528 130170 454598 130226
rect 454654 130170 454722 130226
rect 454778 130170 454848 130226
rect 454528 130102 454848 130170
rect 454528 130046 454598 130102
rect 454654 130046 454722 130102
rect 454778 130046 454848 130102
rect 454528 129978 454848 130046
rect 454528 129922 454598 129978
rect 454654 129922 454722 129978
rect 454778 129922 454848 129978
rect 454528 129888 454848 129922
rect 485248 130350 485568 130384
rect 485248 130294 485318 130350
rect 485374 130294 485442 130350
rect 485498 130294 485568 130350
rect 485248 130226 485568 130294
rect 485248 130170 485318 130226
rect 485374 130170 485442 130226
rect 485498 130170 485568 130226
rect 485248 130102 485568 130170
rect 485248 130046 485318 130102
rect 485374 130046 485442 130102
rect 485498 130046 485568 130102
rect 485248 129978 485568 130046
rect 485248 129922 485318 129978
rect 485374 129922 485442 129978
rect 485498 129922 485568 129978
rect 485248 129888 485568 129922
rect 515968 130350 516288 130384
rect 515968 130294 516038 130350
rect 516094 130294 516162 130350
rect 516218 130294 516288 130350
rect 515968 130226 516288 130294
rect 515968 130170 516038 130226
rect 516094 130170 516162 130226
rect 516218 130170 516288 130226
rect 515968 130102 516288 130170
rect 515968 130046 516038 130102
rect 516094 130046 516162 130102
rect 516218 130046 516288 130102
rect 515968 129978 516288 130046
rect 515968 129922 516038 129978
rect 516094 129922 516162 129978
rect 516218 129922 516288 129978
rect 515968 129888 516288 129922
rect 525154 130350 525774 147922
rect 525154 130294 525250 130350
rect 525306 130294 525374 130350
rect 525430 130294 525498 130350
rect 525554 130294 525622 130350
rect 525678 130294 525774 130350
rect 525154 130226 525774 130294
rect 525154 130170 525250 130226
rect 525306 130170 525374 130226
rect 525430 130170 525498 130226
rect 525554 130170 525622 130226
rect 525678 130170 525774 130226
rect 525154 130102 525774 130170
rect 525154 130046 525250 130102
rect 525306 130046 525374 130102
rect 525430 130046 525498 130102
rect 525554 130046 525622 130102
rect 525678 130046 525774 130102
rect 525154 129978 525774 130046
rect 525154 129922 525250 129978
rect 525306 129922 525374 129978
rect 525430 129922 525498 129978
rect 525554 129922 525622 129978
rect 525678 129922 525774 129978
rect 6874 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 7494 118350
rect 6874 118226 7494 118294
rect 6874 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 7494 118226
rect 6874 118102 7494 118170
rect 6874 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 7494 118102
rect 6874 117978 7494 118046
rect 6874 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 7494 117978
rect 6874 100350 7494 117922
rect 39808 118350 40128 118384
rect 39808 118294 39878 118350
rect 39934 118294 40002 118350
rect 40058 118294 40128 118350
rect 39808 118226 40128 118294
rect 39808 118170 39878 118226
rect 39934 118170 40002 118226
rect 40058 118170 40128 118226
rect 39808 118102 40128 118170
rect 39808 118046 39878 118102
rect 39934 118046 40002 118102
rect 40058 118046 40128 118102
rect 39808 117978 40128 118046
rect 39808 117922 39878 117978
rect 39934 117922 40002 117978
rect 40058 117922 40128 117978
rect 39808 117888 40128 117922
rect 70528 118350 70848 118384
rect 70528 118294 70598 118350
rect 70654 118294 70722 118350
rect 70778 118294 70848 118350
rect 70528 118226 70848 118294
rect 70528 118170 70598 118226
rect 70654 118170 70722 118226
rect 70778 118170 70848 118226
rect 70528 118102 70848 118170
rect 70528 118046 70598 118102
rect 70654 118046 70722 118102
rect 70778 118046 70848 118102
rect 70528 117978 70848 118046
rect 70528 117922 70598 117978
rect 70654 117922 70722 117978
rect 70778 117922 70848 117978
rect 70528 117888 70848 117922
rect 101248 118350 101568 118384
rect 101248 118294 101318 118350
rect 101374 118294 101442 118350
rect 101498 118294 101568 118350
rect 101248 118226 101568 118294
rect 101248 118170 101318 118226
rect 101374 118170 101442 118226
rect 101498 118170 101568 118226
rect 101248 118102 101568 118170
rect 101248 118046 101318 118102
rect 101374 118046 101442 118102
rect 101498 118046 101568 118102
rect 101248 117978 101568 118046
rect 101248 117922 101318 117978
rect 101374 117922 101442 117978
rect 101498 117922 101568 117978
rect 101248 117888 101568 117922
rect 131968 118350 132288 118384
rect 131968 118294 132038 118350
rect 132094 118294 132162 118350
rect 132218 118294 132288 118350
rect 131968 118226 132288 118294
rect 131968 118170 132038 118226
rect 132094 118170 132162 118226
rect 132218 118170 132288 118226
rect 131968 118102 132288 118170
rect 131968 118046 132038 118102
rect 132094 118046 132162 118102
rect 132218 118046 132288 118102
rect 131968 117978 132288 118046
rect 131968 117922 132038 117978
rect 132094 117922 132162 117978
rect 132218 117922 132288 117978
rect 131968 117888 132288 117922
rect 162688 118350 163008 118384
rect 162688 118294 162758 118350
rect 162814 118294 162882 118350
rect 162938 118294 163008 118350
rect 162688 118226 163008 118294
rect 162688 118170 162758 118226
rect 162814 118170 162882 118226
rect 162938 118170 163008 118226
rect 162688 118102 163008 118170
rect 162688 118046 162758 118102
rect 162814 118046 162882 118102
rect 162938 118046 163008 118102
rect 162688 117978 163008 118046
rect 162688 117922 162758 117978
rect 162814 117922 162882 117978
rect 162938 117922 163008 117978
rect 162688 117888 163008 117922
rect 193408 118350 193728 118384
rect 193408 118294 193478 118350
rect 193534 118294 193602 118350
rect 193658 118294 193728 118350
rect 193408 118226 193728 118294
rect 193408 118170 193478 118226
rect 193534 118170 193602 118226
rect 193658 118170 193728 118226
rect 193408 118102 193728 118170
rect 193408 118046 193478 118102
rect 193534 118046 193602 118102
rect 193658 118046 193728 118102
rect 193408 117978 193728 118046
rect 193408 117922 193478 117978
rect 193534 117922 193602 117978
rect 193658 117922 193728 117978
rect 193408 117888 193728 117922
rect 224128 118350 224448 118384
rect 224128 118294 224198 118350
rect 224254 118294 224322 118350
rect 224378 118294 224448 118350
rect 224128 118226 224448 118294
rect 224128 118170 224198 118226
rect 224254 118170 224322 118226
rect 224378 118170 224448 118226
rect 224128 118102 224448 118170
rect 224128 118046 224198 118102
rect 224254 118046 224322 118102
rect 224378 118046 224448 118102
rect 224128 117978 224448 118046
rect 224128 117922 224198 117978
rect 224254 117922 224322 117978
rect 224378 117922 224448 117978
rect 224128 117888 224448 117922
rect 254848 118350 255168 118384
rect 254848 118294 254918 118350
rect 254974 118294 255042 118350
rect 255098 118294 255168 118350
rect 254848 118226 255168 118294
rect 254848 118170 254918 118226
rect 254974 118170 255042 118226
rect 255098 118170 255168 118226
rect 254848 118102 255168 118170
rect 254848 118046 254918 118102
rect 254974 118046 255042 118102
rect 255098 118046 255168 118102
rect 254848 117978 255168 118046
rect 254848 117922 254918 117978
rect 254974 117922 255042 117978
rect 255098 117922 255168 117978
rect 254848 117888 255168 117922
rect 285568 118350 285888 118384
rect 285568 118294 285638 118350
rect 285694 118294 285762 118350
rect 285818 118294 285888 118350
rect 285568 118226 285888 118294
rect 285568 118170 285638 118226
rect 285694 118170 285762 118226
rect 285818 118170 285888 118226
rect 285568 118102 285888 118170
rect 285568 118046 285638 118102
rect 285694 118046 285762 118102
rect 285818 118046 285888 118102
rect 285568 117978 285888 118046
rect 285568 117922 285638 117978
rect 285694 117922 285762 117978
rect 285818 117922 285888 117978
rect 285568 117888 285888 117922
rect 316288 118350 316608 118384
rect 316288 118294 316358 118350
rect 316414 118294 316482 118350
rect 316538 118294 316608 118350
rect 316288 118226 316608 118294
rect 316288 118170 316358 118226
rect 316414 118170 316482 118226
rect 316538 118170 316608 118226
rect 316288 118102 316608 118170
rect 316288 118046 316358 118102
rect 316414 118046 316482 118102
rect 316538 118046 316608 118102
rect 316288 117978 316608 118046
rect 316288 117922 316358 117978
rect 316414 117922 316482 117978
rect 316538 117922 316608 117978
rect 316288 117888 316608 117922
rect 347008 118350 347328 118384
rect 347008 118294 347078 118350
rect 347134 118294 347202 118350
rect 347258 118294 347328 118350
rect 347008 118226 347328 118294
rect 347008 118170 347078 118226
rect 347134 118170 347202 118226
rect 347258 118170 347328 118226
rect 347008 118102 347328 118170
rect 347008 118046 347078 118102
rect 347134 118046 347202 118102
rect 347258 118046 347328 118102
rect 347008 117978 347328 118046
rect 347008 117922 347078 117978
rect 347134 117922 347202 117978
rect 347258 117922 347328 117978
rect 347008 117888 347328 117922
rect 377728 118350 378048 118384
rect 377728 118294 377798 118350
rect 377854 118294 377922 118350
rect 377978 118294 378048 118350
rect 377728 118226 378048 118294
rect 377728 118170 377798 118226
rect 377854 118170 377922 118226
rect 377978 118170 378048 118226
rect 377728 118102 378048 118170
rect 377728 118046 377798 118102
rect 377854 118046 377922 118102
rect 377978 118046 378048 118102
rect 377728 117978 378048 118046
rect 377728 117922 377798 117978
rect 377854 117922 377922 117978
rect 377978 117922 378048 117978
rect 377728 117888 378048 117922
rect 408448 118350 408768 118384
rect 408448 118294 408518 118350
rect 408574 118294 408642 118350
rect 408698 118294 408768 118350
rect 408448 118226 408768 118294
rect 408448 118170 408518 118226
rect 408574 118170 408642 118226
rect 408698 118170 408768 118226
rect 408448 118102 408768 118170
rect 408448 118046 408518 118102
rect 408574 118046 408642 118102
rect 408698 118046 408768 118102
rect 408448 117978 408768 118046
rect 408448 117922 408518 117978
rect 408574 117922 408642 117978
rect 408698 117922 408768 117978
rect 408448 117888 408768 117922
rect 439168 118350 439488 118384
rect 439168 118294 439238 118350
rect 439294 118294 439362 118350
rect 439418 118294 439488 118350
rect 439168 118226 439488 118294
rect 439168 118170 439238 118226
rect 439294 118170 439362 118226
rect 439418 118170 439488 118226
rect 439168 118102 439488 118170
rect 439168 118046 439238 118102
rect 439294 118046 439362 118102
rect 439418 118046 439488 118102
rect 439168 117978 439488 118046
rect 439168 117922 439238 117978
rect 439294 117922 439362 117978
rect 439418 117922 439488 117978
rect 439168 117888 439488 117922
rect 469888 118350 470208 118384
rect 469888 118294 469958 118350
rect 470014 118294 470082 118350
rect 470138 118294 470208 118350
rect 469888 118226 470208 118294
rect 469888 118170 469958 118226
rect 470014 118170 470082 118226
rect 470138 118170 470208 118226
rect 469888 118102 470208 118170
rect 469888 118046 469958 118102
rect 470014 118046 470082 118102
rect 470138 118046 470208 118102
rect 469888 117978 470208 118046
rect 469888 117922 469958 117978
rect 470014 117922 470082 117978
rect 470138 117922 470208 117978
rect 469888 117888 470208 117922
rect 500608 118350 500928 118384
rect 500608 118294 500678 118350
rect 500734 118294 500802 118350
rect 500858 118294 500928 118350
rect 500608 118226 500928 118294
rect 500608 118170 500678 118226
rect 500734 118170 500802 118226
rect 500858 118170 500928 118226
rect 500608 118102 500928 118170
rect 500608 118046 500678 118102
rect 500734 118046 500802 118102
rect 500858 118046 500928 118102
rect 500608 117978 500928 118046
rect 500608 117922 500678 117978
rect 500734 117922 500802 117978
rect 500858 117922 500928 117978
rect 500608 117888 500928 117922
rect 24448 112350 24768 112384
rect 24448 112294 24518 112350
rect 24574 112294 24642 112350
rect 24698 112294 24768 112350
rect 24448 112226 24768 112294
rect 24448 112170 24518 112226
rect 24574 112170 24642 112226
rect 24698 112170 24768 112226
rect 24448 112102 24768 112170
rect 24448 112046 24518 112102
rect 24574 112046 24642 112102
rect 24698 112046 24768 112102
rect 24448 111978 24768 112046
rect 24448 111922 24518 111978
rect 24574 111922 24642 111978
rect 24698 111922 24768 111978
rect 24448 111888 24768 111922
rect 55168 112350 55488 112384
rect 55168 112294 55238 112350
rect 55294 112294 55362 112350
rect 55418 112294 55488 112350
rect 55168 112226 55488 112294
rect 55168 112170 55238 112226
rect 55294 112170 55362 112226
rect 55418 112170 55488 112226
rect 55168 112102 55488 112170
rect 55168 112046 55238 112102
rect 55294 112046 55362 112102
rect 55418 112046 55488 112102
rect 55168 111978 55488 112046
rect 55168 111922 55238 111978
rect 55294 111922 55362 111978
rect 55418 111922 55488 111978
rect 55168 111888 55488 111922
rect 85888 112350 86208 112384
rect 85888 112294 85958 112350
rect 86014 112294 86082 112350
rect 86138 112294 86208 112350
rect 85888 112226 86208 112294
rect 85888 112170 85958 112226
rect 86014 112170 86082 112226
rect 86138 112170 86208 112226
rect 85888 112102 86208 112170
rect 85888 112046 85958 112102
rect 86014 112046 86082 112102
rect 86138 112046 86208 112102
rect 85888 111978 86208 112046
rect 85888 111922 85958 111978
rect 86014 111922 86082 111978
rect 86138 111922 86208 111978
rect 85888 111888 86208 111922
rect 116608 112350 116928 112384
rect 116608 112294 116678 112350
rect 116734 112294 116802 112350
rect 116858 112294 116928 112350
rect 116608 112226 116928 112294
rect 116608 112170 116678 112226
rect 116734 112170 116802 112226
rect 116858 112170 116928 112226
rect 116608 112102 116928 112170
rect 116608 112046 116678 112102
rect 116734 112046 116802 112102
rect 116858 112046 116928 112102
rect 116608 111978 116928 112046
rect 116608 111922 116678 111978
rect 116734 111922 116802 111978
rect 116858 111922 116928 111978
rect 116608 111888 116928 111922
rect 147328 112350 147648 112384
rect 147328 112294 147398 112350
rect 147454 112294 147522 112350
rect 147578 112294 147648 112350
rect 147328 112226 147648 112294
rect 147328 112170 147398 112226
rect 147454 112170 147522 112226
rect 147578 112170 147648 112226
rect 147328 112102 147648 112170
rect 147328 112046 147398 112102
rect 147454 112046 147522 112102
rect 147578 112046 147648 112102
rect 147328 111978 147648 112046
rect 147328 111922 147398 111978
rect 147454 111922 147522 111978
rect 147578 111922 147648 111978
rect 147328 111888 147648 111922
rect 178048 112350 178368 112384
rect 178048 112294 178118 112350
rect 178174 112294 178242 112350
rect 178298 112294 178368 112350
rect 178048 112226 178368 112294
rect 178048 112170 178118 112226
rect 178174 112170 178242 112226
rect 178298 112170 178368 112226
rect 178048 112102 178368 112170
rect 178048 112046 178118 112102
rect 178174 112046 178242 112102
rect 178298 112046 178368 112102
rect 178048 111978 178368 112046
rect 178048 111922 178118 111978
rect 178174 111922 178242 111978
rect 178298 111922 178368 111978
rect 178048 111888 178368 111922
rect 208768 112350 209088 112384
rect 208768 112294 208838 112350
rect 208894 112294 208962 112350
rect 209018 112294 209088 112350
rect 208768 112226 209088 112294
rect 208768 112170 208838 112226
rect 208894 112170 208962 112226
rect 209018 112170 209088 112226
rect 208768 112102 209088 112170
rect 208768 112046 208838 112102
rect 208894 112046 208962 112102
rect 209018 112046 209088 112102
rect 208768 111978 209088 112046
rect 208768 111922 208838 111978
rect 208894 111922 208962 111978
rect 209018 111922 209088 111978
rect 208768 111888 209088 111922
rect 239488 112350 239808 112384
rect 239488 112294 239558 112350
rect 239614 112294 239682 112350
rect 239738 112294 239808 112350
rect 239488 112226 239808 112294
rect 239488 112170 239558 112226
rect 239614 112170 239682 112226
rect 239738 112170 239808 112226
rect 239488 112102 239808 112170
rect 239488 112046 239558 112102
rect 239614 112046 239682 112102
rect 239738 112046 239808 112102
rect 239488 111978 239808 112046
rect 239488 111922 239558 111978
rect 239614 111922 239682 111978
rect 239738 111922 239808 111978
rect 239488 111888 239808 111922
rect 270208 112350 270528 112384
rect 270208 112294 270278 112350
rect 270334 112294 270402 112350
rect 270458 112294 270528 112350
rect 270208 112226 270528 112294
rect 270208 112170 270278 112226
rect 270334 112170 270402 112226
rect 270458 112170 270528 112226
rect 270208 112102 270528 112170
rect 270208 112046 270278 112102
rect 270334 112046 270402 112102
rect 270458 112046 270528 112102
rect 270208 111978 270528 112046
rect 270208 111922 270278 111978
rect 270334 111922 270402 111978
rect 270458 111922 270528 111978
rect 270208 111888 270528 111922
rect 300928 112350 301248 112384
rect 300928 112294 300998 112350
rect 301054 112294 301122 112350
rect 301178 112294 301248 112350
rect 300928 112226 301248 112294
rect 300928 112170 300998 112226
rect 301054 112170 301122 112226
rect 301178 112170 301248 112226
rect 300928 112102 301248 112170
rect 300928 112046 300998 112102
rect 301054 112046 301122 112102
rect 301178 112046 301248 112102
rect 300928 111978 301248 112046
rect 300928 111922 300998 111978
rect 301054 111922 301122 111978
rect 301178 111922 301248 111978
rect 300928 111888 301248 111922
rect 331648 112350 331968 112384
rect 331648 112294 331718 112350
rect 331774 112294 331842 112350
rect 331898 112294 331968 112350
rect 331648 112226 331968 112294
rect 331648 112170 331718 112226
rect 331774 112170 331842 112226
rect 331898 112170 331968 112226
rect 331648 112102 331968 112170
rect 331648 112046 331718 112102
rect 331774 112046 331842 112102
rect 331898 112046 331968 112102
rect 331648 111978 331968 112046
rect 331648 111922 331718 111978
rect 331774 111922 331842 111978
rect 331898 111922 331968 111978
rect 331648 111888 331968 111922
rect 362368 112350 362688 112384
rect 362368 112294 362438 112350
rect 362494 112294 362562 112350
rect 362618 112294 362688 112350
rect 362368 112226 362688 112294
rect 362368 112170 362438 112226
rect 362494 112170 362562 112226
rect 362618 112170 362688 112226
rect 362368 112102 362688 112170
rect 362368 112046 362438 112102
rect 362494 112046 362562 112102
rect 362618 112046 362688 112102
rect 362368 111978 362688 112046
rect 362368 111922 362438 111978
rect 362494 111922 362562 111978
rect 362618 111922 362688 111978
rect 362368 111888 362688 111922
rect 393088 112350 393408 112384
rect 393088 112294 393158 112350
rect 393214 112294 393282 112350
rect 393338 112294 393408 112350
rect 393088 112226 393408 112294
rect 393088 112170 393158 112226
rect 393214 112170 393282 112226
rect 393338 112170 393408 112226
rect 393088 112102 393408 112170
rect 393088 112046 393158 112102
rect 393214 112046 393282 112102
rect 393338 112046 393408 112102
rect 393088 111978 393408 112046
rect 393088 111922 393158 111978
rect 393214 111922 393282 111978
rect 393338 111922 393408 111978
rect 393088 111888 393408 111922
rect 423808 112350 424128 112384
rect 423808 112294 423878 112350
rect 423934 112294 424002 112350
rect 424058 112294 424128 112350
rect 423808 112226 424128 112294
rect 423808 112170 423878 112226
rect 423934 112170 424002 112226
rect 424058 112170 424128 112226
rect 423808 112102 424128 112170
rect 423808 112046 423878 112102
rect 423934 112046 424002 112102
rect 424058 112046 424128 112102
rect 423808 111978 424128 112046
rect 423808 111922 423878 111978
rect 423934 111922 424002 111978
rect 424058 111922 424128 111978
rect 423808 111888 424128 111922
rect 454528 112350 454848 112384
rect 454528 112294 454598 112350
rect 454654 112294 454722 112350
rect 454778 112294 454848 112350
rect 454528 112226 454848 112294
rect 454528 112170 454598 112226
rect 454654 112170 454722 112226
rect 454778 112170 454848 112226
rect 454528 112102 454848 112170
rect 454528 112046 454598 112102
rect 454654 112046 454722 112102
rect 454778 112046 454848 112102
rect 454528 111978 454848 112046
rect 454528 111922 454598 111978
rect 454654 111922 454722 111978
rect 454778 111922 454848 111978
rect 454528 111888 454848 111922
rect 485248 112350 485568 112384
rect 485248 112294 485318 112350
rect 485374 112294 485442 112350
rect 485498 112294 485568 112350
rect 485248 112226 485568 112294
rect 485248 112170 485318 112226
rect 485374 112170 485442 112226
rect 485498 112170 485568 112226
rect 485248 112102 485568 112170
rect 485248 112046 485318 112102
rect 485374 112046 485442 112102
rect 485498 112046 485568 112102
rect 485248 111978 485568 112046
rect 485248 111922 485318 111978
rect 485374 111922 485442 111978
rect 485498 111922 485568 111978
rect 485248 111888 485568 111922
rect 515968 112350 516288 112384
rect 515968 112294 516038 112350
rect 516094 112294 516162 112350
rect 516218 112294 516288 112350
rect 515968 112226 516288 112294
rect 515968 112170 516038 112226
rect 516094 112170 516162 112226
rect 516218 112170 516288 112226
rect 515968 112102 516288 112170
rect 515968 112046 516038 112102
rect 516094 112046 516162 112102
rect 516218 112046 516288 112102
rect 515968 111978 516288 112046
rect 515968 111922 516038 111978
rect 516094 111922 516162 111978
rect 516218 111922 516288 111978
rect 515968 111888 516288 111922
rect 525154 112350 525774 129922
rect 525154 112294 525250 112350
rect 525306 112294 525374 112350
rect 525430 112294 525498 112350
rect 525554 112294 525622 112350
rect 525678 112294 525774 112350
rect 525154 112226 525774 112294
rect 525154 112170 525250 112226
rect 525306 112170 525374 112226
rect 525430 112170 525498 112226
rect 525554 112170 525622 112226
rect 525678 112170 525774 112226
rect 525154 112102 525774 112170
rect 525154 112046 525250 112102
rect 525306 112046 525374 112102
rect 525430 112046 525498 112102
rect 525554 112046 525622 112102
rect 525678 112046 525774 112102
rect 525154 111978 525774 112046
rect 525154 111922 525250 111978
rect 525306 111922 525374 111978
rect 525430 111922 525498 111978
rect 525554 111922 525622 111978
rect 525678 111922 525774 111978
rect 6874 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 7494 100350
rect 6874 100226 7494 100294
rect 6874 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 7494 100226
rect 6874 100102 7494 100170
rect 6874 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 7494 100102
rect 6874 99978 7494 100046
rect 6874 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 7494 99978
rect 6874 82350 7494 99922
rect 39808 100350 40128 100384
rect 39808 100294 39878 100350
rect 39934 100294 40002 100350
rect 40058 100294 40128 100350
rect 39808 100226 40128 100294
rect 39808 100170 39878 100226
rect 39934 100170 40002 100226
rect 40058 100170 40128 100226
rect 39808 100102 40128 100170
rect 39808 100046 39878 100102
rect 39934 100046 40002 100102
rect 40058 100046 40128 100102
rect 39808 99978 40128 100046
rect 39808 99922 39878 99978
rect 39934 99922 40002 99978
rect 40058 99922 40128 99978
rect 39808 99888 40128 99922
rect 70528 100350 70848 100384
rect 70528 100294 70598 100350
rect 70654 100294 70722 100350
rect 70778 100294 70848 100350
rect 70528 100226 70848 100294
rect 70528 100170 70598 100226
rect 70654 100170 70722 100226
rect 70778 100170 70848 100226
rect 70528 100102 70848 100170
rect 70528 100046 70598 100102
rect 70654 100046 70722 100102
rect 70778 100046 70848 100102
rect 70528 99978 70848 100046
rect 70528 99922 70598 99978
rect 70654 99922 70722 99978
rect 70778 99922 70848 99978
rect 70528 99888 70848 99922
rect 101248 100350 101568 100384
rect 101248 100294 101318 100350
rect 101374 100294 101442 100350
rect 101498 100294 101568 100350
rect 101248 100226 101568 100294
rect 101248 100170 101318 100226
rect 101374 100170 101442 100226
rect 101498 100170 101568 100226
rect 101248 100102 101568 100170
rect 101248 100046 101318 100102
rect 101374 100046 101442 100102
rect 101498 100046 101568 100102
rect 101248 99978 101568 100046
rect 101248 99922 101318 99978
rect 101374 99922 101442 99978
rect 101498 99922 101568 99978
rect 101248 99888 101568 99922
rect 131968 100350 132288 100384
rect 131968 100294 132038 100350
rect 132094 100294 132162 100350
rect 132218 100294 132288 100350
rect 131968 100226 132288 100294
rect 131968 100170 132038 100226
rect 132094 100170 132162 100226
rect 132218 100170 132288 100226
rect 131968 100102 132288 100170
rect 131968 100046 132038 100102
rect 132094 100046 132162 100102
rect 132218 100046 132288 100102
rect 131968 99978 132288 100046
rect 131968 99922 132038 99978
rect 132094 99922 132162 99978
rect 132218 99922 132288 99978
rect 131968 99888 132288 99922
rect 162688 100350 163008 100384
rect 162688 100294 162758 100350
rect 162814 100294 162882 100350
rect 162938 100294 163008 100350
rect 162688 100226 163008 100294
rect 162688 100170 162758 100226
rect 162814 100170 162882 100226
rect 162938 100170 163008 100226
rect 162688 100102 163008 100170
rect 162688 100046 162758 100102
rect 162814 100046 162882 100102
rect 162938 100046 163008 100102
rect 162688 99978 163008 100046
rect 162688 99922 162758 99978
rect 162814 99922 162882 99978
rect 162938 99922 163008 99978
rect 162688 99888 163008 99922
rect 193408 100350 193728 100384
rect 193408 100294 193478 100350
rect 193534 100294 193602 100350
rect 193658 100294 193728 100350
rect 193408 100226 193728 100294
rect 193408 100170 193478 100226
rect 193534 100170 193602 100226
rect 193658 100170 193728 100226
rect 193408 100102 193728 100170
rect 193408 100046 193478 100102
rect 193534 100046 193602 100102
rect 193658 100046 193728 100102
rect 193408 99978 193728 100046
rect 193408 99922 193478 99978
rect 193534 99922 193602 99978
rect 193658 99922 193728 99978
rect 193408 99888 193728 99922
rect 224128 100350 224448 100384
rect 224128 100294 224198 100350
rect 224254 100294 224322 100350
rect 224378 100294 224448 100350
rect 224128 100226 224448 100294
rect 224128 100170 224198 100226
rect 224254 100170 224322 100226
rect 224378 100170 224448 100226
rect 224128 100102 224448 100170
rect 224128 100046 224198 100102
rect 224254 100046 224322 100102
rect 224378 100046 224448 100102
rect 224128 99978 224448 100046
rect 224128 99922 224198 99978
rect 224254 99922 224322 99978
rect 224378 99922 224448 99978
rect 224128 99888 224448 99922
rect 254848 100350 255168 100384
rect 254848 100294 254918 100350
rect 254974 100294 255042 100350
rect 255098 100294 255168 100350
rect 254848 100226 255168 100294
rect 254848 100170 254918 100226
rect 254974 100170 255042 100226
rect 255098 100170 255168 100226
rect 254848 100102 255168 100170
rect 254848 100046 254918 100102
rect 254974 100046 255042 100102
rect 255098 100046 255168 100102
rect 254848 99978 255168 100046
rect 254848 99922 254918 99978
rect 254974 99922 255042 99978
rect 255098 99922 255168 99978
rect 254848 99888 255168 99922
rect 285568 100350 285888 100384
rect 285568 100294 285638 100350
rect 285694 100294 285762 100350
rect 285818 100294 285888 100350
rect 285568 100226 285888 100294
rect 285568 100170 285638 100226
rect 285694 100170 285762 100226
rect 285818 100170 285888 100226
rect 285568 100102 285888 100170
rect 285568 100046 285638 100102
rect 285694 100046 285762 100102
rect 285818 100046 285888 100102
rect 285568 99978 285888 100046
rect 285568 99922 285638 99978
rect 285694 99922 285762 99978
rect 285818 99922 285888 99978
rect 285568 99888 285888 99922
rect 316288 100350 316608 100384
rect 316288 100294 316358 100350
rect 316414 100294 316482 100350
rect 316538 100294 316608 100350
rect 316288 100226 316608 100294
rect 316288 100170 316358 100226
rect 316414 100170 316482 100226
rect 316538 100170 316608 100226
rect 316288 100102 316608 100170
rect 316288 100046 316358 100102
rect 316414 100046 316482 100102
rect 316538 100046 316608 100102
rect 316288 99978 316608 100046
rect 316288 99922 316358 99978
rect 316414 99922 316482 99978
rect 316538 99922 316608 99978
rect 316288 99888 316608 99922
rect 347008 100350 347328 100384
rect 347008 100294 347078 100350
rect 347134 100294 347202 100350
rect 347258 100294 347328 100350
rect 347008 100226 347328 100294
rect 347008 100170 347078 100226
rect 347134 100170 347202 100226
rect 347258 100170 347328 100226
rect 347008 100102 347328 100170
rect 347008 100046 347078 100102
rect 347134 100046 347202 100102
rect 347258 100046 347328 100102
rect 347008 99978 347328 100046
rect 347008 99922 347078 99978
rect 347134 99922 347202 99978
rect 347258 99922 347328 99978
rect 347008 99888 347328 99922
rect 377728 100350 378048 100384
rect 377728 100294 377798 100350
rect 377854 100294 377922 100350
rect 377978 100294 378048 100350
rect 377728 100226 378048 100294
rect 377728 100170 377798 100226
rect 377854 100170 377922 100226
rect 377978 100170 378048 100226
rect 377728 100102 378048 100170
rect 377728 100046 377798 100102
rect 377854 100046 377922 100102
rect 377978 100046 378048 100102
rect 377728 99978 378048 100046
rect 377728 99922 377798 99978
rect 377854 99922 377922 99978
rect 377978 99922 378048 99978
rect 377728 99888 378048 99922
rect 408448 100350 408768 100384
rect 408448 100294 408518 100350
rect 408574 100294 408642 100350
rect 408698 100294 408768 100350
rect 408448 100226 408768 100294
rect 408448 100170 408518 100226
rect 408574 100170 408642 100226
rect 408698 100170 408768 100226
rect 408448 100102 408768 100170
rect 408448 100046 408518 100102
rect 408574 100046 408642 100102
rect 408698 100046 408768 100102
rect 408448 99978 408768 100046
rect 408448 99922 408518 99978
rect 408574 99922 408642 99978
rect 408698 99922 408768 99978
rect 408448 99888 408768 99922
rect 439168 100350 439488 100384
rect 439168 100294 439238 100350
rect 439294 100294 439362 100350
rect 439418 100294 439488 100350
rect 439168 100226 439488 100294
rect 439168 100170 439238 100226
rect 439294 100170 439362 100226
rect 439418 100170 439488 100226
rect 439168 100102 439488 100170
rect 439168 100046 439238 100102
rect 439294 100046 439362 100102
rect 439418 100046 439488 100102
rect 439168 99978 439488 100046
rect 439168 99922 439238 99978
rect 439294 99922 439362 99978
rect 439418 99922 439488 99978
rect 439168 99888 439488 99922
rect 469888 100350 470208 100384
rect 469888 100294 469958 100350
rect 470014 100294 470082 100350
rect 470138 100294 470208 100350
rect 469888 100226 470208 100294
rect 469888 100170 469958 100226
rect 470014 100170 470082 100226
rect 470138 100170 470208 100226
rect 469888 100102 470208 100170
rect 469888 100046 469958 100102
rect 470014 100046 470082 100102
rect 470138 100046 470208 100102
rect 469888 99978 470208 100046
rect 469888 99922 469958 99978
rect 470014 99922 470082 99978
rect 470138 99922 470208 99978
rect 469888 99888 470208 99922
rect 500608 100350 500928 100384
rect 500608 100294 500678 100350
rect 500734 100294 500802 100350
rect 500858 100294 500928 100350
rect 500608 100226 500928 100294
rect 500608 100170 500678 100226
rect 500734 100170 500802 100226
rect 500858 100170 500928 100226
rect 500608 100102 500928 100170
rect 500608 100046 500678 100102
rect 500734 100046 500802 100102
rect 500858 100046 500928 100102
rect 500608 99978 500928 100046
rect 500608 99922 500678 99978
rect 500734 99922 500802 99978
rect 500858 99922 500928 99978
rect 500608 99888 500928 99922
rect 24448 94350 24768 94384
rect 24448 94294 24518 94350
rect 24574 94294 24642 94350
rect 24698 94294 24768 94350
rect 24448 94226 24768 94294
rect 24448 94170 24518 94226
rect 24574 94170 24642 94226
rect 24698 94170 24768 94226
rect 24448 94102 24768 94170
rect 24448 94046 24518 94102
rect 24574 94046 24642 94102
rect 24698 94046 24768 94102
rect 24448 93978 24768 94046
rect 24448 93922 24518 93978
rect 24574 93922 24642 93978
rect 24698 93922 24768 93978
rect 24448 93888 24768 93922
rect 55168 94350 55488 94384
rect 55168 94294 55238 94350
rect 55294 94294 55362 94350
rect 55418 94294 55488 94350
rect 55168 94226 55488 94294
rect 55168 94170 55238 94226
rect 55294 94170 55362 94226
rect 55418 94170 55488 94226
rect 55168 94102 55488 94170
rect 55168 94046 55238 94102
rect 55294 94046 55362 94102
rect 55418 94046 55488 94102
rect 55168 93978 55488 94046
rect 55168 93922 55238 93978
rect 55294 93922 55362 93978
rect 55418 93922 55488 93978
rect 55168 93888 55488 93922
rect 85888 94350 86208 94384
rect 85888 94294 85958 94350
rect 86014 94294 86082 94350
rect 86138 94294 86208 94350
rect 85888 94226 86208 94294
rect 85888 94170 85958 94226
rect 86014 94170 86082 94226
rect 86138 94170 86208 94226
rect 85888 94102 86208 94170
rect 85888 94046 85958 94102
rect 86014 94046 86082 94102
rect 86138 94046 86208 94102
rect 85888 93978 86208 94046
rect 85888 93922 85958 93978
rect 86014 93922 86082 93978
rect 86138 93922 86208 93978
rect 85888 93888 86208 93922
rect 116608 94350 116928 94384
rect 116608 94294 116678 94350
rect 116734 94294 116802 94350
rect 116858 94294 116928 94350
rect 116608 94226 116928 94294
rect 116608 94170 116678 94226
rect 116734 94170 116802 94226
rect 116858 94170 116928 94226
rect 116608 94102 116928 94170
rect 116608 94046 116678 94102
rect 116734 94046 116802 94102
rect 116858 94046 116928 94102
rect 116608 93978 116928 94046
rect 116608 93922 116678 93978
rect 116734 93922 116802 93978
rect 116858 93922 116928 93978
rect 116608 93888 116928 93922
rect 147328 94350 147648 94384
rect 147328 94294 147398 94350
rect 147454 94294 147522 94350
rect 147578 94294 147648 94350
rect 147328 94226 147648 94294
rect 147328 94170 147398 94226
rect 147454 94170 147522 94226
rect 147578 94170 147648 94226
rect 147328 94102 147648 94170
rect 147328 94046 147398 94102
rect 147454 94046 147522 94102
rect 147578 94046 147648 94102
rect 147328 93978 147648 94046
rect 147328 93922 147398 93978
rect 147454 93922 147522 93978
rect 147578 93922 147648 93978
rect 147328 93888 147648 93922
rect 178048 94350 178368 94384
rect 178048 94294 178118 94350
rect 178174 94294 178242 94350
rect 178298 94294 178368 94350
rect 178048 94226 178368 94294
rect 178048 94170 178118 94226
rect 178174 94170 178242 94226
rect 178298 94170 178368 94226
rect 178048 94102 178368 94170
rect 178048 94046 178118 94102
rect 178174 94046 178242 94102
rect 178298 94046 178368 94102
rect 178048 93978 178368 94046
rect 178048 93922 178118 93978
rect 178174 93922 178242 93978
rect 178298 93922 178368 93978
rect 178048 93888 178368 93922
rect 208768 94350 209088 94384
rect 208768 94294 208838 94350
rect 208894 94294 208962 94350
rect 209018 94294 209088 94350
rect 208768 94226 209088 94294
rect 208768 94170 208838 94226
rect 208894 94170 208962 94226
rect 209018 94170 209088 94226
rect 208768 94102 209088 94170
rect 208768 94046 208838 94102
rect 208894 94046 208962 94102
rect 209018 94046 209088 94102
rect 208768 93978 209088 94046
rect 208768 93922 208838 93978
rect 208894 93922 208962 93978
rect 209018 93922 209088 93978
rect 208768 93888 209088 93922
rect 239488 94350 239808 94384
rect 239488 94294 239558 94350
rect 239614 94294 239682 94350
rect 239738 94294 239808 94350
rect 239488 94226 239808 94294
rect 239488 94170 239558 94226
rect 239614 94170 239682 94226
rect 239738 94170 239808 94226
rect 239488 94102 239808 94170
rect 239488 94046 239558 94102
rect 239614 94046 239682 94102
rect 239738 94046 239808 94102
rect 239488 93978 239808 94046
rect 239488 93922 239558 93978
rect 239614 93922 239682 93978
rect 239738 93922 239808 93978
rect 239488 93888 239808 93922
rect 270208 94350 270528 94384
rect 270208 94294 270278 94350
rect 270334 94294 270402 94350
rect 270458 94294 270528 94350
rect 270208 94226 270528 94294
rect 270208 94170 270278 94226
rect 270334 94170 270402 94226
rect 270458 94170 270528 94226
rect 270208 94102 270528 94170
rect 270208 94046 270278 94102
rect 270334 94046 270402 94102
rect 270458 94046 270528 94102
rect 270208 93978 270528 94046
rect 270208 93922 270278 93978
rect 270334 93922 270402 93978
rect 270458 93922 270528 93978
rect 270208 93888 270528 93922
rect 300928 94350 301248 94384
rect 300928 94294 300998 94350
rect 301054 94294 301122 94350
rect 301178 94294 301248 94350
rect 300928 94226 301248 94294
rect 300928 94170 300998 94226
rect 301054 94170 301122 94226
rect 301178 94170 301248 94226
rect 300928 94102 301248 94170
rect 300928 94046 300998 94102
rect 301054 94046 301122 94102
rect 301178 94046 301248 94102
rect 300928 93978 301248 94046
rect 300928 93922 300998 93978
rect 301054 93922 301122 93978
rect 301178 93922 301248 93978
rect 300928 93888 301248 93922
rect 331648 94350 331968 94384
rect 331648 94294 331718 94350
rect 331774 94294 331842 94350
rect 331898 94294 331968 94350
rect 331648 94226 331968 94294
rect 331648 94170 331718 94226
rect 331774 94170 331842 94226
rect 331898 94170 331968 94226
rect 331648 94102 331968 94170
rect 331648 94046 331718 94102
rect 331774 94046 331842 94102
rect 331898 94046 331968 94102
rect 331648 93978 331968 94046
rect 331648 93922 331718 93978
rect 331774 93922 331842 93978
rect 331898 93922 331968 93978
rect 331648 93888 331968 93922
rect 362368 94350 362688 94384
rect 362368 94294 362438 94350
rect 362494 94294 362562 94350
rect 362618 94294 362688 94350
rect 362368 94226 362688 94294
rect 362368 94170 362438 94226
rect 362494 94170 362562 94226
rect 362618 94170 362688 94226
rect 362368 94102 362688 94170
rect 362368 94046 362438 94102
rect 362494 94046 362562 94102
rect 362618 94046 362688 94102
rect 362368 93978 362688 94046
rect 362368 93922 362438 93978
rect 362494 93922 362562 93978
rect 362618 93922 362688 93978
rect 362368 93888 362688 93922
rect 393088 94350 393408 94384
rect 393088 94294 393158 94350
rect 393214 94294 393282 94350
rect 393338 94294 393408 94350
rect 393088 94226 393408 94294
rect 393088 94170 393158 94226
rect 393214 94170 393282 94226
rect 393338 94170 393408 94226
rect 393088 94102 393408 94170
rect 393088 94046 393158 94102
rect 393214 94046 393282 94102
rect 393338 94046 393408 94102
rect 393088 93978 393408 94046
rect 393088 93922 393158 93978
rect 393214 93922 393282 93978
rect 393338 93922 393408 93978
rect 393088 93888 393408 93922
rect 423808 94350 424128 94384
rect 423808 94294 423878 94350
rect 423934 94294 424002 94350
rect 424058 94294 424128 94350
rect 423808 94226 424128 94294
rect 423808 94170 423878 94226
rect 423934 94170 424002 94226
rect 424058 94170 424128 94226
rect 423808 94102 424128 94170
rect 423808 94046 423878 94102
rect 423934 94046 424002 94102
rect 424058 94046 424128 94102
rect 423808 93978 424128 94046
rect 423808 93922 423878 93978
rect 423934 93922 424002 93978
rect 424058 93922 424128 93978
rect 423808 93888 424128 93922
rect 454528 94350 454848 94384
rect 454528 94294 454598 94350
rect 454654 94294 454722 94350
rect 454778 94294 454848 94350
rect 454528 94226 454848 94294
rect 454528 94170 454598 94226
rect 454654 94170 454722 94226
rect 454778 94170 454848 94226
rect 454528 94102 454848 94170
rect 454528 94046 454598 94102
rect 454654 94046 454722 94102
rect 454778 94046 454848 94102
rect 454528 93978 454848 94046
rect 454528 93922 454598 93978
rect 454654 93922 454722 93978
rect 454778 93922 454848 93978
rect 454528 93888 454848 93922
rect 485248 94350 485568 94384
rect 485248 94294 485318 94350
rect 485374 94294 485442 94350
rect 485498 94294 485568 94350
rect 485248 94226 485568 94294
rect 485248 94170 485318 94226
rect 485374 94170 485442 94226
rect 485498 94170 485568 94226
rect 485248 94102 485568 94170
rect 485248 94046 485318 94102
rect 485374 94046 485442 94102
rect 485498 94046 485568 94102
rect 485248 93978 485568 94046
rect 485248 93922 485318 93978
rect 485374 93922 485442 93978
rect 485498 93922 485568 93978
rect 485248 93888 485568 93922
rect 515968 94350 516288 94384
rect 515968 94294 516038 94350
rect 516094 94294 516162 94350
rect 516218 94294 516288 94350
rect 515968 94226 516288 94294
rect 515968 94170 516038 94226
rect 516094 94170 516162 94226
rect 516218 94170 516288 94226
rect 515968 94102 516288 94170
rect 515968 94046 516038 94102
rect 516094 94046 516162 94102
rect 516218 94046 516288 94102
rect 515968 93978 516288 94046
rect 515968 93922 516038 93978
rect 516094 93922 516162 93978
rect 516218 93922 516288 93978
rect 515968 93888 516288 93922
rect 525154 94350 525774 111922
rect 525154 94294 525250 94350
rect 525306 94294 525374 94350
rect 525430 94294 525498 94350
rect 525554 94294 525622 94350
rect 525678 94294 525774 94350
rect 525154 94226 525774 94294
rect 525154 94170 525250 94226
rect 525306 94170 525374 94226
rect 525430 94170 525498 94226
rect 525554 94170 525622 94226
rect 525678 94170 525774 94226
rect 525154 94102 525774 94170
rect 525154 94046 525250 94102
rect 525306 94046 525374 94102
rect 525430 94046 525498 94102
rect 525554 94046 525622 94102
rect 525678 94046 525774 94102
rect 525154 93978 525774 94046
rect 525154 93922 525250 93978
rect 525306 93922 525374 93978
rect 525430 93922 525498 93978
rect 525554 93922 525622 93978
rect 525678 93922 525774 93978
rect 6874 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 7494 82350
rect 6874 82226 7494 82294
rect 6874 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 7494 82226
rect 6874 82102 7494 82170
rect 6874 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 7494 82102
rect 6874 81978 7494 82046
rect 6874 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 7494 81978
rect 6874 64350 7494 81922
rect 39808 82350 40128 82384
rect 39808 82294 39878 82350
rect 39934 82294 40002 82350
rect 40058 82294 40128 82350
rect 39808 82226 40128 82294
rect 39808 82170 39878 82226
rect 39934 82170 40002 82226
rect 40058 82170 40128 82226
rect 39808 82102 40128 82170
rect 39808 82046 39878 82102
rect 39934 82046 40002 82102
rect 40058 82046 40128 82102
rect 39808 81978 40128 82046
rect 39808 81922 39878 81978
rect 39934 81922 40002 81978
rect 40058 81922 40128 81978
rect 39808 81888 40128 81922
rect 70528 82350 70848 82384
rect 70528 82294 70598 82350
rect 70654 82294 70722 82350
rect 70778 82294 70848 82350
rect 70528 82226 70848 82294
rect 70528 82170 70598 82226
rect 70654 82170 70722 82226
rect 70778 82170 70848 82226
rect 70528 82102 70848 82170
rect 70528 82046 70598 82102
rect 70654 82046 70722 82102
rect 70778 82046 70848 82102
rect 70528 81978 70848 82046
rect 70528 81922 70598 81978
rect 70654 81922 70722 81978
rect 70778 81922 70848 81978
rect 70528 81888 70848 81922
rect 101248 82350 101568 82384
rect 101248 82294 101318 82350
rect 101374 82294 101442 82350
rect 101498 82294 101568 82350
rect 101248 82226 101568 82294
rect 101248 82170 101318 82226
rect 101374 82170 101442 82226
rect 101498 82170 101568 82226
rect 101248 82102 101568 82170
rect 101248 82046 101318 82102
rect 101374 82046 101442 82102
rect 101498 82046 101568 82102
rect 101248 81978 101568 82046
rect 101248 81922 101318 81978
rect 101374 81922 101442 81978
rect 101498 81922 101568 81978
rect 101248 81888 101568 81922
rect 131968 82350 132288 82384
rect 131968 82294 132038 82350
rect 132094 82294 132162 82350
rect 132218 82294 132288 82350
rect 131968 82226 132288 82294
rect 131968 82170 132038 82226
rect 132094 82170 132162 82226
rect 132218 82170 132288 82226
rect 131968 82102 132288 82170
rect 131968 82046 132038 82102
rect 132094 82046 132162 82102
rect 132218 82046 132288 82102
rect 131968 81978 132288 82046
rect 131968 81922 132038 81978
rect 132094 81922 132162 81978
rect 132218 81922 132288 81978
rect 131968 81888 132288 81922
rect 162688 82350 163008 82384
rect 162688 82294 162758 82350
rect 162814 82294 162882 82350
rect 162938 82294 163008 82350
rect 162688 82226 163008 82294
rect 162688 82170 162758 82226
rect 162814 82170 162882 82226
rect 162938 82170 163008 82226
rect 162688 82102 163008 82170
rect 162688 82046 162758 82102
rect 162814 82046 162882 82102
rect 162938 82046 163008 82102
rect 162688 81978 163008 82046
rect 162688 81922 162758 81978
rect 162814 81922 162882 81978
rect 162938 81922 163008 81978
rect 162688 81888 163008 81922
rect 193408 82350 193728 82384
rect 193408 82294 193478 82350
rect 193534 82294 193602 82350
rect 193658 82294 193728 82350
rect 193408 82226 193728 82294
rect 193408 82170 193478 82226
rect 193534 82170 193602 82226
rect 193658 82170 193728 82226
rect 193408 82102 193728 82170
rect 193408 82046 193478 82102
rect 193534 82046 193602 82102
rect 193658 82046 193728 82102
rect 193408 81978 193728 82046
rect 193408 81922 193478 81978
rect 193534 81922 193602 81978
rect 193658 81922 193728 81978
rect 193408 81888 193728 81922
rect 224128 82350 224448 82384
rect 224128 82294 224198 82350
rect 224254 82294 224322 82350
rect 224378 82294 224448 82350
rect 224128 82226 224448 82294
rect 224128 82170 224198 82226
rect 224254 82170 224322 82226
rect 224378 82170 224448 82226
rect 224128 82102 224448 82170
rect 224128 82046 224198 82102
rect 224254 82046 224322 82102
rect 224378 82046 224448 82102
rect 224128 81978 224448 82046
rect 224128 81922 224198 81978
rect 224254 81922 224322 81978
rect 224378 81922 224448 81978
rect 224128 81888 224448 81922
rect 254848 82350 255168 82384
rect 254848 82294 254918 82350
rect 254974 82294 255042 82350
rect 255098 82294 255168 82350
rect 254848 82226 255168 82294
rect 254848 82170 254918 82226
rect 254974 82170 255042 82226
rect 255098 82170 255168 82226
rect 254848 82102 255168 82170
rect 254848 82046 254918 82102
rect 254974 82046 255042 82102
rect 255098 82046 255168 82102
rect 254848 81978 255168 82046
rect 254848 81922 254918 81978
rect 254974 81922 255042 81978
rect 255098 81922 255168 81978
rect 254848 81888 255168 81922
rect 285568 82350 285888 82384
rect 285568 82294 285638 82350
rect 285694 82294 285762 82350
rect 285818 82294 285888 82350
rect 285568 82226 285888 82294
rect 285568 82170 285638 82226
rect 285694 82170 285762 82226
rect 285818 82170 285888 82226
rect 285568 82102 285888 82170
rect 285568 82046 285638 82102
rect 285694 82046 285762 82102
rect 285818 82046 285888 82102
rect 285568 81978 285888 82046
rect 285568 81922 285638 81978
rect 285694 81922 285762 81978
rect 285818 81922 285888 81978
rect 285568 81888 285888 81922
rect 316288 82350 316608 82384
rect 316288 82294 316358 82350
rect 316414 82294 316482 82350
rect 316538 82294 316608 82350
rect 316288 82226 316608 82294
rect 316288 82170 316358 82226
rect 316414 82170 316482 82226
rect 316538 82170 316608 82226
rect 316288 82102 316608 82170
rect 316288 82046 316358 82102
rect 316414 82046 316482 82102
rect 316538 82046 316608 82102
rect 316288 81978 316608 82046
rect 316288 81922 316358 81978
rect 316414 81922 316482 81978
rect 316538 81922 316608 81978
rect 316288 81888 316608 81922
rect 347008 82350 347328 82384
rect 347008 82294 347078 82350
rect 347134 82294 347202 82350
rect 347258 82294 347328 82350
rect 347008 82226 347328 82294
rect 347008 82170 347078 82226
rect 347134 82170 347202 82226
rect 347258 82170 347328 82226
rect 347008 82102 347328 82170
rect 347008 82046 347078 82102
rect 347134 82046 347202 82102
rect 347258 82046 347328 82102
rect 347008 81978 347328 82046
rect 347008 81922 347078 81978
rect 347134 81922 347202 81978
rect 347258 81922 347328 81978
rect 347008 81888 347328 81922
rect 377728 82350 378048 82384
rect 377728 82294 377798 82350
rect 377854 82294 377922 82350
rect 377978 82294 378048 82350
rect 377728 82226 378048 82294
rect 377728 82170 377798 82226
rect 377854 82170 377922 82226
rect 377978 82170 378048 82226
rect 377728 82102 378048 82170
rect 377728 82046 377798 82102
rect 377854 82046 377922 82102
rect 377978 82046 378048 82102
rect 377728 81978 378048 82046
rect 377728 81922 377798 81978
rect 377854 81922 377922 81978
rect 377978 81922 378048 81978
rect 377728 81888 378048 81922
rect 408448 82350 408768 82384
rect 408448 82294 408518 82350
rect 408574 82294 408642 82350
rect 408698 82294 408768 82350
rect 408448 82226 408768 82294
rect 408448 82170 408518 82226
rect 408574 82170 408642 82226
rect 408698 82170 408768 82226
rect 408448 82102 408768 82170
rect 408448 82046 408518 82102
rect 408574 82046 408642 82102
rect 408698 82046 408768 82102
rect 408448 81978 408768 82046
rect 408448 81922 408518 81978
rect 408574 81922 408642 81978
rect 408698 81922 408768 81978
rect 408448 81888 408768 81922
rect 439168 82350 439488 82384
rect 439168 82294 439238 82350
rect 439294 82294 439362 82350
rect 439418 82294 439488 82350
rect 439168 82226 439488 82294
rect 439168 82170 439238 82226
rect 439294 82170 439362 82226
rect 439418 82170 439488 82226
rect 439168 82102 439488 82170
rect 439168 82046 439238 82102
rect 439294 82046 439362 82102
rect 439418 82046 439488 82102
rect 439168 81978 439488 82046
rect 439168 81922 439238 81978
rect 439294 81922 439362 81978
rect 439418 81922 439488 81978
rect 439168 81888 439488 81922
rect 469888 82350 470208 82384
rect 469888 82294 469958 82350
rect 470014 82294 470082 82350
rect 470138 82294 470208 82350
rect 469888 82226 470208 82294
rect 469888 82170 469958 82226
rect 470014 82170 470082 82226
rect 470138 82170 470208 82226
rect 469888 82102 470208 82170
rect 469888 82046 469958 82102
rect 470014 82046 470082 82102
rect 470138 82046 470208 82102
rect 469888 81978 470208 82046
rect 469888 81922 469958 81978
rect 470014 81922 470082 81978
rect 470138 81922 470208 81978
rect 469888 81888 470208 81922
rect 500608 82350 500928 82384
rect 500608 82294 500678 82350
rect 500734 82294 500802 82350
rect 500858 82294 500928 82350
rect 500608 82226 500928 82294
rect 500608 82170 500678 82226
rect 500734 82170 500802 82226
rect 500858 82170 500928 82226
rect 500608 82102 500928 82170
rect 500608 82046 500678 82102
rect 500734 82046 500802 82102
rect 500858 82046 500928 82102
rect 500608 81978 500928 82046
rect 500608 81922 500678 81978
rect 500734 81922 500802 81978
rect 500858 81922 500928 81978
rect 500608 81888 500928 81922
rect 24448 76350 24768 76384
rect 24448 76294 24518 76350
rect 24574 76294 24642 76350
rect 24698 76294 24768 76350
rect 24448 76226 24768 76294
rect 24448 76170 24518 76226
rect 24574 76170 24642 76226
rect 24698 76170 24768 76226
rect 24448 76102 24768 76170
rect 24448 76046 24518 76102
rect 24574 76046 24642 76102
rect 24698 76046 24768 76102
rect 24448 75978 24768 76046
rect 24448 75922 24518 75978
rect 24574 75922 24642 75978
rect 24698 75922 24768 75978
rect 24448 75888 24768 75922
rect 55168 76350 55488 76384
rect 55168 76294 55238 76350
rect 55294 76294 55362 76350
rect 55418 76294 55488 76350
rect 55168 76226 55488 76294
rect 55168 76170 55238 76226
rect 55294 76170 55362 76226
rect 55418 76170 55488 76226
rect 55168 76102 55488 76170
rect 55168 76046 55238 76102
rect 55294 76046 55362 76102
rect 55418 76046 55488 76102
rect 55168 75978 55488 76046
rect 55168 75922 55238 75978
rect 55294 75922 55362 75978
rect 55418 75922 55488 75978
rect 55168 75888 55488 75922
rect 85888 76350 86208 76384
rect 85888 76294 85958 76350
rect 86014 76294 86082 76350
rect 86138 76294 86208 76350
rect 85888 76226 86208 76294
rect 85888 76170 85958 76226
rect 86014 76170 86082 76226
rect 86138 76170 86208 76226
rect 85888 76102 86208 76170
rect 85888 76046 85958 76102
rect 86014 76046 86082 76102
rect 86138 76046 86208 76102
rect 85888 75978 86208 76046
rect 85888 75922 85958 75978
rect 86014 75922 86082 75978
rect 86138 75922 86208 75978
rect 85888 75888 86208 75922
rect 116608 76350 116928 76384
rect 116608 76294 116678 76350
rect 116734 76294 116802 76350
rect 116858 76294 116928 76350
rect 116608 76226 116928 76294
rect 116608 76170 116678 76226
rect 116734 76170 116802 76226
rect 116858 76170 116928 76226
rect 116608 76102 116928 76170
rect 116608 76046 116678 76102
rect 116734 76046 116802 76102
rect 116858 76046 116928 76102
rect 116608 75978 116928 76046
rect 116608 75922 116678 75978
rect 116734 75922 116802 75978
rect 116858 75922 116928 75978
rect 116608 75888 116928 75922
rect 147328 76350 147648 76384
rect 147328 76294 147398 76350
rect 147454 76294 147522 76350
rect 147578 76294 147648 76350
rect 147328 76226 147648 76294
rect 147328 76170 147398 76226
rect 147454 76170 147522 76226
rect 147578 76170 147648 76226
rect 147328 76102 147648 76170
rect 147328 76046 147398 76102
rect 147454 76046 147522 76102
rect 147578 76046 147648 76102
rect 147328 75978 147648 76046
rect 147328 75922 147398 75978
rect 147454 75922 147522 75978
rect 147578 75922 147648 75978
rect 147328 75888 147648 75922
rect 178048 76350 178368 76384
rect 178048 76294 178118 76350
rect 178174 76294 178242 76350
rect 178298 76294 178368 76350
rect 178048 76226 178368 76294
rect 178048 76170 178118 76226
rect 178174 76170 178242 76226
rect 178298 76170 178368 76226
rect 178048 76102 178368 76170
rect 178048 76046 178118 76102
rect 178174 76046 178242 76102
rect 178298 76046 178368 76102
rect 178048 75978 178368 76046
rect 178048 75922 178118 75978
rect 178174 75922 178242 75978
rect 178298 75922 178368 75978
rect 178048 75888 178368 75922
rect 208768 76350 209088 76384
rect 208768 76294 208838 76350
rect 208894 76294 208962 76350
rect 209018 76294 209088 76350
rect 208768 76226 209088 76294
rect 208768 76170 208838 76226
rect 208894 76170 208962 76226
rect 209018 76170 209088 76226
rect 208768 76102 209088 76170
rect 208768 76046 208838 76102
rect 208894 76046 208962 76102
rect 209018 76046 209088 76102
rect 208768 75978 209088 76046
rect 208768 75922 208838 75978
rect 208894 75922 208962 75978
rect 209018 75922 209088 75978
rect 208768 75888 209088 75922
rect 239488 76350 239808 76384
rect 239488 76294 239558 76350
rect 239614 76294 239682 76350
rect 239738 76294 239808 76350
rect 239488 76226 239808 76294
rect 239488 76170 239558 76226
rect 239614 76170 239682 76226
rect 239738 76170 239808 76226
rect 239488 76102 239808 76170
rect 239488 76046 239558 76102
rect 239614 76046 239682 76102
rect 239738 76046 239808 76102
rect 239488 75978 239808 76046
rect 239488 75922 239558 75978
rect 239614 75922 239682 75978
rect 239738 75922 239808 75978
rect 239488 75888 239808 75922
rect 270208 76350 270528 76384
rect 270208 76294 270278 76350
rect 270334 76294 270402 76350
rect 270458 76294 270528 76350
rect 270208 76226 270528 76294
rect 270208 76170 270278 76226
rect 270334 76170 270402 76226
rect 270458 76170 270528 76226
rect 270208 76102 270528 76170
rect 270208 76046 270278 76102
rect 270334 76046 270402 76102
rect 270458 76046 270528 76102
rect 270208 75978 270528 76046
rect 270208 75922 270278 75978
rect 270334 75922 270402 75978
rect 270458 75922 270528 75978
rect 270208 75888 270528 75922
rect 300928 76350 301248 76384
rect 300928 76294 300998 76350
rect 301054 76294 301122 76350
rect 301178 76294 301248 76350
rect 300928 76226 301248 76294
rect 300928 76170 300998 76226
rect 301054 76170 301122 76226
rect 301178 76170 301248 76226
rect 300928 76102 301248 76170
rect 300928 76046 300998 76102
rect 301054 76046 301122 76102
rect 301178 76046 301248 76102
rect 300928 75978 301248 76046
rect 300928 75922 300998 75978
rect 301054 75922 301122 75978
rect 301178 75922 301248 75978
rect 300928 75888 301248 75922
rect 331648 76350 331968 76384
rect 331648 76294 331718 76350
rect 331774 76294 331842 76350
rect 331898 76294 331968 76350
rect 331648 76226 331968 76294
rect 331648 76170 331718 76226
rect 331774 76170 331842 76226
rect 331898 76170 331968 76226
rect 331648 76102 331968 76170
rect 331648 76046 331718 76102
rect 331774 76046 331842 76102
rect 331898 76046 331968 76102
rect 331648 75978 331968 76046
rect 331648 75922 331718 75978
rect 331774 75922 331842 75978
rect 331898 75922 331968 75978
rect 331648 75888 331968 75922
rect 362368 76350 362688 76384
rect 362368 76294 362438 76350
rect 362494 76294 362562 76350
rect 362618 76294 362688 76350
rect 362368 76226 362688 76294
rect 362368 76170 362438 76226
rect 362494 76170 362562 76226
rect 362618 76170 362688 76226
rect 362368 76102 362688 76170
rect 362368 76046 362438 76102
rect 362494 76046 362562 76102
rect 362618 76046 362688 76102
rect 362368 75978 362688 76046
rect 362368 75922 362438 75978
rect 362494 75922 362562 75978
rect 362618 75922 362688 75978
rect 362368 75888 362688 75922
rect 393088 76350 393408 76384
rect 393088 76294 393158 76350
rect 393214 76294 393282 76350
rect 393338 76294 393408 76350
rect 393088 76226 393408 76294
rect 393088 76170 393158 76226
rect 393214 76170 393282 76226
rect 393338 76170 393408 76226
rect 393088 76102 393408 76170
rect 393088 76046 393158 76102
rect 393214 76046 393282 76102
rect 393338 76046 393408 76102
rect 393088 75978 393408 76046
rect 393088 75922 393158 75978
rect 393214 75922 393282 75978
rect 393338 75922 393408 75978
rect 393088 75888 393408 75922
rect 423808 76350 424128 76384
rect 423808 76294 423878 76350
rect 423934 76294 424002 76350
rect 424058 76294 424128 76350
rect 423808 76226 424128 76294
rect 423808 76170 423878 76226
rect 423934 76170 424002 76226
rect 424058 76170 424128 76226
rect 423808 76102 424128 76170
rect 423808 76046 423878 76102
rect 423934 76046 424002 76102
rect 424058 76046 424128 76102
rect 423808 75978 424128 76046
rect 423808 75922 423878 75978
rect 423934 75922 424002 75978
rect 424058 75922 424128 75978
rect 423808 75888 424128 75922
rect 454528 76350 454848 76384
rect 454528 76294 454598 76350
rect 454654 76294 454722 76350
rect 454778 76294 454848 76350
rect 454528 76226 454848 76294
rect 454528 76170 454598 76226
rect 454654 76170 454722 76226
rect 454778 76170 454848 76226
rect 454528 76102 454848 76170
rect 454528 76046 454598 76102
rect 454654 76046 454722 76102
rect 454778 76046 454848 76102
rect 454528 75978 454848 76046
rect 454528 75922 454598 75978
rect 454654 75922 454722 75978
rect 454778 75922 454848 75978
rect 454528 75888 454848 75922
rect 485248 76350 485568 76384
rect 485248 76294 485318 76350
rect 485374 76294 485442 76350
rect 485498 76294 485568 76350
rect 485248 76226 485568 76294
rect 485248 76170 485318 76226
rect 485374 76170 485442 76226
rect 485498 76170 485568 76226
rect 485248 76102 485568 76170
rect 485248 76046 485318 76102
rect 485374 76046 485442 76102
rect 485498 76046 485568 76102
rect 485248 75978 485568 76046
rect 485248 75922 485318 75978
rect 485374 75922 485442 75978
rect 485498 75922 485568 75978
rect 485248 75888 485568 75922
rect 515968 76350 516288 76384
rect 515968 76294 516038 76350
rect 516094 76294 516162 76350
rect 516218 76294 516288 76350
rect 515968 76226 516288 76294
rect 515968 76170 516038 76226
rect 516094 76170 516162 76226
rect 516218 76170 516288 76226
rect 515968 76102 516288 76170
rect 515968 76046 516038 76102
rect 516094 76046 516162 76102
rect 516218 76046 516288 76102
rect 515968 75978 516288 76046
rect 515968 75922 516038 75978
rect 516094 75922 516162 75978
rect 516218 75922 516288 75978
rect 515968 75888 516288 75922
rect 525154 76350 525774 93922
rect 525154 76294 525250 76350
rect 525306 76294 525374 76350
rect 525430 76294 525498 76350
rect 525554 76294 525622 76350
rect 525678 76294 525774 76350
rect 525154 76226 525774 76294
rect 525154 76170 525250 76226
rect 525306 76170 525374 76226
rect 525430 76170 525498 76226
rect 525554 76170 525622 76226
rect 525678 76170 525774 76226
rect 525154 76102 525774 76170
rect 525154 76046 525250 76102
rect 525306 76046 525374 76102
rect 525430 76046 525498 76102
rect 525554 76046 525622 76102
rect 525678 76046 525774 76102
rect 525154 75978 525774 76046
rect 525154 75922 525250 75978
rect 525306 75922 525374 75978
rect 525430 75922 525498 75978
rect 525554 75922 525622 75978
rect 525678 75922 525774 75978
rect 6874 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 7494 64350
rect 6874 64226 7494 64294
rect 6874 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 7494 64226
rect 6874 64102 7494 64170
rect 6874 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 7494 64102
rect 6874 63978 7494 64046
rect 6874 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 7494 63978
rect 6874 46350 7494 63922
rect 39808 64350 40128 64384
rect 39808 64294 39878 64350
rect 39934 64294 40002 64350
rect 40058 64294 40128 64350
rect 39808 64226 40128 64294
rect 39808 64170 39878 64226
rect 39934 64170 40002 64226
rect 40058 64170 40128 64226
rect 39808 64102 40128 64170
rect 39808 64046 39878 64102
rect 39934 64046 40002 64102
rect 40058 64046 40128 64102
rect 39808 63978 40128 64046
rect 39808 63922 39878 63978
rect 39934 63922 40002 63978
rect 40058 63922 40128 63978
rect 39808 63888 40128 63922
rect 70528 64350 70848 64384
rect 70528 64294 70598 64350
rect 70654 64294 70722 64350
rect 70778 64294 70848 64350
rect 70528 64226 70848 64294
rect 70528 64170 70598 64226
rect 70654 64170 70722 64226
rect 70778 64170 70848 64226
rect 70528 64102 70848 64170
rect 70528 64046 70598 64102
rect 70654 64046 70722 64102
rect 70778 64046 70848 64102
rect 70528 63978 70848 64046
rect 70528 63922 70598 63978
rect 70654 63922 70722 63978
rect 70778 63922 70848 63978
rect 70528 63888 70848 63922
rect 101248 64350 101568 64384
rect 101248 64294 101318 64350
rect 101374 64294 101442 64350
rect 101498 64294 101568 64350
rect 101248 64226 101568 64294
rect 101248 64170 101318 64226
rect 101374 64170 101442 64226
rect 101498 64170 101568 64226
rect 101248 64102 101568 64170
rect 101248 64046 101318 64102
rect 101374 64046 101442 64102
rect 101498 64046 101568 64102
rect 101248 63978 101568 64046
rect 101248 63922 101318 63978
rect 101374 63922 101442 63978
rect 101498 63922 101568 63978
rect 101248 63888 101568 63922
rect 131968 64350 132288 64384
rect 131968 64294 132038 64350
rect 132094 64294 132162 64350
rect 132218 64294 132288 64350
rect 131968 64226 132288 64294
rect 131968 64170 132038 64226
rect 132094 64170 132162 64226
rect 132218 64170 132288 64226
rect 131968 64102 132288 64170
rect 131968 64046 132038 64102
rect 132094 64046 132162 64102
rect 132218 64046 132288 64102
rect 131968 63978 132288 64046
rect 131968 63922 132038 63978
rect 132094 63922 132162 63978
rect 132218 63922 132288 63978
rect 131968 63888 132288 63922
rect 162688 64350 163008 64384
rect 162688 64294 162758 64350
rect 162814 64294 162882 64350
rect 162938 64294 163008 64350
rect 162688 64226 163008 64294
rect 162688 64170 162758 64226
rect 162814 64170 162882 64226
rect 162938 64170 163008 64226
rect 162688 64102 163008 64170
rect 162688 64046 162758 64102
rect 162814 64046 162882 64102
rect 162938 64046 163008 64102
rect 162688 63978 163008 64046
rect 162688 63922 162758 63978
rect 162814 63922 162882 63978
rect 162938 63922 163008 63978
rect 162688 63888 163008 63922
rect 193408 64350 193728 64384
rect 193408 64294 193478 64350
rect 193534 64294 193602 64350
rect 193658 64294 193728 64350
rect 193408 64226 193728 64294
rect 193408 64170 193478 64226
rect 193534 64170 193602 64226
rect 193658 64170 193728 64226
rect 193408 64102 193728 64170
rect 193408 64046 193478 64102
rect 193534 64046 193602 64102
rect 193658 64046 193728 64102
rect 193408 63978 193728 64046
rect 193408 63922 193478 63978
rect 193534 63922 193602 63978
rect 193658 63922 193728 63978
rect 193408 63888 193728 63922
rect 224128 64350 224448 64384
rect 224128 64294 224198 64350
rect 224254 64294 224322 64350
rect 224378 64294 224448 64350
rect 224128 64226 224448 64294
rect 224128 64170 224198 64226
rect 224254 64170 224322 64226
rect 224378 64170 224448 64226
rect 224128 64102 224448 64170
rect 224128 64046 224198 64102
rect 224254 64046 224322 64102
rect 224378 64046 224448 64102
rect 224128 63978 224448 64046
rect 224128 63922 224198 63978
rect 224254 63922 224322 63978
rect 224378 63922 224448 63978
rect 224128 63888 224448 63922
rect 254848 64350 255168 64384
rect 254848 64294 254918 64350
rect 254974 64294 255042 64350
rect 255098 64294 255168 64350
rect 254848 64226 255168 64294
rect 254848 64170 254918 64226
rect 254974 64170 255042 64226
rect 255098 64170 255168 64226
rect 254848 64102 255168 64170
rect 254848 64046 254918 64102
rect 254974 64046 255042 64102
rect 255098 64046 255168 64102
rect 254848 63978 255168 64046
rect 254848 63922 254918 63978
rect 254974 63922 255042 63978
rect 255098 63922 255168 63978
rect 254848 63888 255168 63922
rect 285568 64350 285888 64384
rect 285568 64294 285638 64350
rect 285694 64294 285762 64350
rect 285818 64294 285888 64350
rect 285568 64226 285888 64294
rect 285568 64170 285638 64226
rect 285694 64170 285762 64226
rect 285818 64170 285888 64226
rect 285568 64102 285888 64170
rect 285568 64046 285638 64102
rect 285694 64046 285762 64102
rect 285818 64046 285888 64102
rect 285568 63978 285888 64046
rect 285568 63922 285638 63978
rect 285694 63922 285762 63978
rect 285818 63922 285888 63978
rect 285568 63888 285888 63922
rect 316288 64350 316608 64384
rect 316288 64294 316358 64350
rect 316414 64294 316482 64350
rect 316538 64294 316608 64350
rect 316288 64226 316608 64294
rect 316288 64170 316358 64226
rect 316414 64170 316482 64226
rect 316538 64170 316608 64226
rect 316288 64102 316608 64170
rect 316288 64046 316358 64102
rect 316414 64046 316482 64102
rect 316538 64046 316608 64102
rect 316288 63978 316608 64046
rect 316288 63922 316358 63978
rect 316414 63922 316482 63978
rect 316538 63922 316608 63978
rect 316288 63888 316608 63922
rect 347008 64350 347328 64384
rect 347008 64294 347078 64350
rect 347134 64294 347202 64350
rect 347258 64294 347328 64350
rect 347008 64226 347328 64294
rect 347008 64170 347078 64226
rect 347134 64170 347202 64226
rect 347258 64170 347328 64226
rect 347008 64102 347328 64170
rect 347008 64046 347078 64102
rect 347134 64046 347202 64102
rect 347258 64046 347328 64102
rect 347008 63978 347328 64046
rect 347008 63922 347078 63978
rect 347134 63922 347202 63978
rect 347258 63922 347328 63978
rect 347008 63888 347328 63922
rect 377728 64350 378048 64384
rect 377728 64294 377798 64350
rect 377854 64294 377922 64350
rect 377978 64294 378048 64350
rect 377728 64226 378048 64294
rect 377728 64170 377798 64226
rect 377854 64170 377922 64226
rect 377978 64170 378048 64226
rect 377728 64102 378048 64170
rect 377728 64046 377798 64102
rect 377854 64046 377922 64102
rect 377978 64046 378048 64102
rect 377728 63978 378048 64046
rect 377728 63922 377798 63978
rect 377854 63922 377922 63978
rect 377978 63922 378048 63978
rect 377728 63888 378048 63922
rect 408448 64350 408768 64384
rect 408448 64294 408518 64350
rect 408574 64294 408642 64350
rect 408698 64294 408768 64350
rect 408448 64226 408768 64294
rect 408448 64170 408518 64226
rect 408574 64170 408642 64226
rect 408698 64170 408768 64226
rect 408448 64102 408768 64170
rect 408448 64046 408518 64102
rect 408574 64046 408642 64102
rect 408698 64046 408768 64102
rect 408448 63978 408768 64046
rect 408448 63922 408518 63978
rect 408574 63922 408642 63978
rect 408698 63922 408768 63978
rect 408448 63888 408768 63922
rect 439168 64350 439488 64384
rect 439168 64294 439238 64350
rect 439294 64294 439362 64350
rect 439418 64294 439488 64350
rect 439168 64226 439488 64294
rect 439168 64170 439238 64226
rect 439294 64170 439362 64226
rect 439418 64170 439488 64226
rect 439168 64102 439488 64170
rect 439168 64046 439238 64102
rect 439294 64046 439362 64102
rect 439418 64046 439488 64102
rect 439168 63978 439488 64046
rect 439168 63922 439238 63978
rect 439294 63922 439362 63978
rect 439418 63922 439488 63978
rect 439168 63888 439488 63922
rect 469888 64350 470208 64384
rect 469888 64294 469958 64350
rect 470014 64294 470082 64350
rect 470138 64294 470208 64350
rect 469888 64226 470208 64294
rect 469888 64170 469958 64226
rect 470014 64170 470082 64226
rect 470138 64170 470208 64226
rect 469888 64102 470208 64170
rect 469888 64046 469958 64102
rect 470014 64046 470082 64102
rect 470138 64046 470208 64102
rect 469888 63978 470208 64046
rect 469888 63922 469958 63978
rect 470014 63922 470082 63978
rect 470138 63922 470208 63978
rect 469888 63888 470208 63922
rect 500608 64350 500928 64384
rect 500608 64294 500678 64350
rect 500734 64294 500802 64350
rect 500858 64294 500928 64350
rect 500608 64226 500928 64294
rect 500608 64170 500678 64226
rect 500734 64170 500802 64226
rect 500858 64170 500928 64226
rect 500608 64102 500928 64170
rect 500608 64046 500678 64102
rect 500734 64046 500802 64102
rect 500858 64046 500928 64102
rect 500608 63978 500928 64046
rect 500608 63922 500678 63978
rect 500734 63922 500802 63978
rect 500858 63922 500928 63978
rect 500608 63888 500928 63922
rect 24448 58350 24768 58384
rect 24448 58294 24518 58350
rect 24574 58294 24642 58350
rect 24698 58294 24768 58350
rect 24448 58226 24768 58294
rect 24448 58170 24518 58226
rect 24574 58170 24642 58226
rect 24698 58170 24768 58226
rect 24448 58102 24768 58170
rect 24448 58046 24518 58102
rect 24574 58046 24642 58102
rect 24698 58046 24768 58102
rect 24448 57978 24768 58046
rect 24448 57922 24518 57978
rect 24574 57922 24642 57978
rect 24698 57922 24768 57978
rect 24448 57888 24768 57922
rect 55168 58350 55488 58384
rect 55168 58294 55238 58350
rect 55294 58294 55362 58350
rect 55418 58294 55488 58350
rect 55168 58226 55488 58294
rect 55168 58170 55238 58226
rect 55294 58170 55362 58226
rect 55418 58170 55488 58226
rect 55168 58102 55488 58170
rect 55168 58046 55238 58102
rect 55294 58046 55362 58102
rect 55418 58046 55488 58102
rect 55168 57978 55488 58046
rect 55168 57922 55238 57978
rect 55294 57922 55362 57978
rect 55418 57922 55488 57978
rect 55168 57888 55488 57922
rect 85888 58350 86208 58384
rect 85888 58294 85958 58350
rect 86014 58294 86082 58350
rect 86138 58294 86208 58350
rect 85888 58226 86208 58294
rect 85888 58170 85958 58226
rect 86014 58170 86082 58226
rect 86138 58170 86208 58226
rect 85888 58102 86208 58170
rect 85888 58046 85958 58102
rect 86014 58046 86082 58102
rect 86138 58046 86208 58102
rect 85888 57978 86208 58046
rect 85888 57922 85958 57978
rect 86014 57922 86082 57978
rect 86138 57922 86208 57978
rect 85888 57888 86208 57922
rect 116608 58350 116928 58384
rect 116608 58294 116678 58350
rect 116734 58294 116802 58350
rect 116858 58294 116928 58350
rect 116608 58226 116928 58294
rect 116608 58170 116678 58226
rect 116734 58170 116802 58226
rect 116858 58170 116928 58226
rect 116608 58102 116928 58170
rect 116608 58046 116678 58102
rect 116734 58046 116802 58102
rect 116858 58046 116928 58102
rect 116608 57978 116928 58046
rect 116608 57922 116678 57978
rect 116734 57922 116802 57978
rect 116858 57922 116928 57978
rect 116608 57888 116928 57922
rect 147328 58350 147648 58384
rect 147328 58294 147398 58350
rect 147454 58294 147522 58350
rect 147578 58294 147648 58350
rect 147328 58226 147648 58294
rect 147328 58170 147398 58226
rect 147454 58170 147522 58226
rect 147578 58170 147648 58226
rect 147328 58102 147648 58170
rect 147328 58046 147398 58102
rect 147454 58046 147522 58102
rect 147578 58046 147648 58102
rect 147328 57978 147648 58046
rect 147328 57922 147398 57978
rect 147454 57922 147522 57978
rect 147578 57922 147648 57978
rect 147328 57888 147648 57922
rect 178048 58350 178368 58384
rect 178048 58294 178118 58350
rect 178174 58294 178242 58350
rect 178298 58294 178368 58350
rect 178048 58226 178368 58294
rect 178048 58170 178118 58226
rect 178174 58170 178242 58226
rect 178298 58170 178368 58226
rect 178048 58102 178368 58170
rect 178048 58046 178118 58102
rect 178174 58046 178242 58102
rect 178298 58046 178368 58102
rect 178048 57978 178368 58046
rect 178048 57922 178118 57978
rect 178174 57922 178242 57978
rect 178298 57922 178368 57978
rect 178048 57888 178368 57922
rect 208768 58350 209088 58384
rect 208768 58294 208838 58350
rect 208894 58294 208962 58350
rect 209018 58294 209088 58350
rect 208768 58226 209088 58294
rect 208768 58170 208838 58226
rect 208894 58170 208962 58226
rect 209018 58170 209088 58226
rect 208768 58102 209088 58170
rect 208768 58046 208838 58102
rect 208894 58046 208962 58102
rect 209018 58046 209088 58102
rect 208768 57978 209088 58046
rect 208768 57922 208838 57978
rect 208894 57922 208962 57978
rect 209018 57922 209088 57978
rect 208768 57888 209088 57922
rect 239488 58350 239808 58384
rect 239488 58294 239558 58350
rect 239614 58294 239682 58350
rect 239738 58294 239808 58350
rect 239488 58226 239808 58294
rect 239488 58170 239558 58226
rect 239614 58170 239682 58226
rect 239738 58170 239808 58226
rect 239488 58102 239808 58170
rect 239488 58046 239558 58102
rect 239614 58046 239682 58102
rect 239738 58046 239808 58102
rect 239488 57978 239808 58046
rect 239488 57922 239558 57978
rect 239614 57922 239682 57978
rect 239738 57922 239808 57978
rect 239488 57888 239808 57922
rect 270208 58350 270528 58384
rect 270208 58294 270278 58350
rect 270334 58294 270402 58350
rect 270458 58294 270528 58350
rect 270208 58226 270528 58294
rect 270208 58170 270278 58226
rect 270334 58170 270402 58226
rect 270458 58170 270528 58226
rect 270208 58102 270528 58170
rect 270208 58046 270278 58102
rect 270334 58046 270402 58102
rect 270458 58046 270528 58102
rect 270208 57978 270528 58046
rect 270208 57922 270278 57978
rect 270334 57922 270402 57978
rect 270458 57922 270528 57978
rect 270208 57888 270528 57922
rect 300928 58350 301248 58384
rect 300928 58294 300998 58350
rect 301054 58294 301122 58350
rect 301178 58294 301248 58350
rect 300928 58226 301248 58294
rect 300928 58170 300998 58226
rect 301054 58170 301122 58226
rect 301178 58170 301248 58226
rect 300928 58102 301248 58170
rect 300928 58046 300998 58102
rect 301054 58046 301122 58102
rect 301178 58046 301248 58102
rect 300928 57978 301248 58046
rect 300928 57922 300998 57978
rect 301054 57922 301122 57978
rect 301178 57922 301248 57978
rect 300928 57888 301248 57922
rect 331648 58350 331968 58384
rect 331648 58294 331718 58350
rect 331774 58294 331842 58350
rect 331898 58294 331968 58350
rect 331648 58226 331968 58294
rect 331648 58170 331718 58226
rect 331774 58170 331842 58226
rect 331898 58170 331968 58226
rect 331648 58102 331968 58170
rect 331648 58046 331718 58102
rect 331774 58046 331842 58102
rect 331898 58046 331968 58102
rect 331648 57978 331968 58046
rect 331648 57922 331718 57978
rect 331774 57922 331842 57978
rect 331898 57922 331968 57978
rect 331648 57888 331968 57922
rect 362368 58350 362688 58384
rect 362368 58294 362438 58350
rect 362494 58294 362562 58350
rect 362618 58294 362688 58350
rect 362368 58226 362688 58294
rect 362368 58170 362438 58226
rect 362494 58170 362562 58226
rect 362618 58170 362688 58226
rect 362368 58102 362688 58170
rect 362368 58046 362438 58102
rect 362494 58046 362562 58102
rect 362618 58046 362688 58102
rect 362368 57978 362688 58046
rect 362368 57922 362438 57978
rect 362494 57922 362562 57978
rect 362618 57922 362688 57978
rect 362368 57888 362688 57922
rect 393088 58350 393408 58384
rect 393088 58294 393158 58350
rect 393214 58294 393282 58350
rect 393338 58294 393408 58350
rect 393088 58226 393408 58294
rect 393088 58170 393158 58226
rect 393214 58170 393282 58226
rect 393338 58170 393408 58226
rect 393088 58102 393408 58170
rect 393088 58046 393158 58102
rect 393214 58046 393282 58102
rect 393338 58046 393408 58102
rect 393088 57978 393408 58046
rect 393088 57922 393158 57978
rect 393214 57922 393282 57978
rect 393338 57922 393408 57978
rect 393088 57888 393408 57922
rect 423808 58350 424128 58384
rect 423808 58294 423878 58350
rect 423934 58294 424002 58350
rect 424058 58294 424128 58350
rect 423808 58226 424128 58294
rect 423808 58170 423878 58226
rect 423934 58170 424002 58226
rect 424058 58170 424128 58226
rect 423808 58102 424128 58170
rect 423808 58046 423878 58102
rect 423934 58046 424002 58102
rect 424058 58046 424128 58102
rect 423808 57978 424128 58046
rect 423808 57922 423878 57978
rect 423934 57922 424002 57978
rect 424058 57922 424128 57978
rect 423808 57888 424128 57922
rect 454528 58350 454848 58384
rect 454528 58294 454598 58350
rect 454654 58294 454722 58350
rect 454778 58294 454848 58350
rect 454528 58226 454848 58294
rect 454528 58170 454598 58226
rect 454654 58170 454722 58226
rect 454778 58170 454848 58226
rect 454528 58102 454848 58170
rect 454528 58046 454598 58102
rect 454654 58046 454722 58102
rect 454778 58046 454848 58102
rect 454528 57978 454848 58046
rect 454528 57922 454598 57978
rect 454654 57922 454722 57978
rect 454778 57922 454848 57978
rect 454528 57888 454848 57922
rect 485248 58350 485568 58384
rect 485248 58294 485318 58350
rect 485374 58294 485442 58350
rect 485498 58294 485568 58350
rect 485248 58226 485568 58294
rect 485248 58170 485318 58226
rect 485374 58170 485442 58226
rect 485498 58170 485568 58226
rect 485248 58102 485568 58170
rect 485248 58046 485318 58102
rect 485374 58046 485442 58102
rect 485498 58046 485568 58102
rect 485248 57978 485568 58046
rect 485248 57922 485318 57978
rect 485374 57922 485442 57978
rect 485498 57922 485568 57978
rect 485248 57888 485568 57922
rect 515968 58350 516288 58384
rect 515968 58294 516038 58350
rect 516094 58294 516162 58350
rect 516218 58294 516288 58350
rect 515968 58226 516288 58294
rect 515968 58170 516038 58226
rect 516094 58170 516162 58226
rect 516218 58170 516288 58226
rect 515968 58102 516288 58170
rect 515968 58046 516038 58102
rect 516094 58046 516162 58102
rect 516218 58046 516288 58102
rect 515968 57978 516288 58046
rect 515968 57922 516038 57978
rect 516094 57922 516162 57978
rect 516218 57922 516288 57978
rect 515968 57888 516288 57922
rect 525154 58350 525774 75922
rect 525154 58294 525250 58350
rect 525306 58294 525374 58350
rect 525430 58294 525498 58350
rect 525554 58294 525622 58350
rect 525678 58294 525774 58350
rect 525154 58226 525774 58294
rect 525154 58170 525250 58226
rect 525306 58170 525374 58226
rect 525430 58170 525498 58226
rect 525554 58170 525622 58226
rect 525678 58170 525774 58226
rect 525154 58102 525774 58170
rect 525154 58046 525250 58102
rect 525306 58046 525374 58102
rect 525430 58046 525498 58102
rect 525554 58046 525622 58102
rect 525678 58046 525774 58102
rect 525154 57978 525774 58046
rect 525154 57922 525250 57978
rect 525306 57922 525374 57978
rect 525430 57922 525498 57978
rect 525554 57922 525622 57978
rect 525678 57922 525774 57978
rect 6874 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 7494 46350
rect 6874 46226 7494 46294
rect 6874 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 7494 46226
rect 6874 46102 7494 46170
rect 6874 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 7494 46102
rect 6874 45978 7494 46046
rect 6874 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 7494 45978
rect 6874 28350 7494 45922
rect 39808 46350 40128 46384
rect 39808 46294 39878 46350
rect 39934 46294 40002 46350
rect 40058 46294 40128 46350
rect 39808 46226 40128 46294
rect 39808 46170 39878 46226
rect 39934 46170 40002 46226
rect 40058 46170 40128 46226
rect 39808 46102 40128 46170
rect 39808 46046 39878 46102
rect 39934 46046 40002 46102
rect 40058 46046 40128 46102
rect 39808 45978 40128 46046
rect 39808 45922 39878 45978
rect 39934 45922 40002 45978
rect 40058 45922 40128 45978
rect 39808 45888 40128 45922
rect 70528 46350 70848 46384
rect 70528 46294 70598 46350
rect 70654 46294 70722 46350
rect 70778 46294 70848 46350
rect 70528 46226 70848 46294
rect 70528 46170 70598 46226
rect 70654 46170 70722 46226
rect 70778 46170 70848 46226
rect 70528 46102 70848 46170
rect 70528 46046 70598 46102
rect 70654 46046 70722 46102
rect 70778 46046 70848 46102
rect 70528 45978 70848 46046
rect 70528 45922 70598 45978
rect 70654 45922 70722 45978
rect 70778 45922 70848 45978
rect 70528 45888 70848 45922
rect 101248 46350 101568 46384
rect 101248 46294 101318 46350
rect 101374 46294 101442 46350
rect 101498 46294 101568 46350
rect 101248 46226 101568 46294
rect 101248 46170 101318 46226
rect 101374 46170 101442 46226
rect 101498 46170 101568 46226
rect 101248 46102 101568 46170
rect 101248 46046 101318 46102
rect 101374 46046 101442 46102
rect 101498 46046 101568 46102
rect 101248 45978 101568 46046
rect 101248 45922 101318 45978
rect 101374 45922 101442 45978
rect 101498 45922 101568 45978
rect 101248 45888 101568 45922
rect 131968 46350 132288 46384
rect 131968 46294 132038 46350
rect 132094 46294 132162 46350
rect 132218 46294 132288 46350
rect 131968 46226 132288 46294
rect 131968 46170 132038 46226
rect 132094 46170 132162 46226
rect 132218 46170 132288 46226
rect 131968 46102 132288 46170
rect 131968 46046 132038 46102
rect 132094 46046 132162 46102
rect 132218 46046 132288 46102
rect 131968 45978 132288 46046
rect 131968 45922 132038 45978
rect 132094 45922 132162 45978
rect 132218 45922 132288 45978
rect 131968 45888 132288 45922
rect 162688 46350 163008 46384
rect 162688 46294 162758 46350
rect 162814 46294 162882 46350
rect 162938 46294 163008 46350
rect 162688 46226 163008 46294
rect 162688 46170 162758 46226
rect 162814 46170 162882 46226
rect 162938 46170 163008 46226
rect 162688 46102 163008 46170
rect 162688 46046 162758 46102
rect 162814 46046 162882 46102
rect 162938 46046 163008 46102
rect 162688 45978 163008 46046
rect 162688 45922 162758 45978
rect 162814 45922 162882 45978
rect 162938 45922 163008 45978
rect 162688 45888 163008 45922
rect 193408 46350 193728 46384
rect 193408 46294 193478 46350
rect 193534 46294 193602 46350
rect 193658 46294 193728 46350
rect 193408 46226 193728 46294
rect 193408 46170 193478 46226
rect 193534 46170 193602 46226
rect 193658 46170 193728 46226
rect 193408 46102 193728 46170
rect 193408 46046 193478 46102
rect 193534 46046 193602 46102
rect 193658 46046 193728 46102
rect 193408 45978 193728 46046
rect 193408 45922 193478 45978
rect 193534 45922 193602 45978
rect 193658 45922 193728 45978
rect 193408 45888 193728 45922
rect 224128 46350 224448 46384
rect 224128 46294 224198 46350
rect 224254 46294 224322 46350
rect 224378 46294 224448 46350
rect 224128 46226 224448 46294
rect 224128 46170 224198 46226
rect 224254 46170 224322 46226
rect 224378 46170 224448 46226
rect 224128 46102 224448 46170
rect 224128 46046 224198 46102
rect 224254 46046 224322 46102
rect 224378 46046 224448 46102
rect 224128 45978 224448 46046
rect 224128 45922 224198 45978
rect 224254 45922 224322 45978
rect 224378 45922 224448 45978
rect 224128 45888 224448 45922
rect 254848 46350 255168 46384
rect 254848 46294 254918 46350
rect 254974 46294 255042 46350
rect 255098 46294 255168 46350
rect 254848 46226 255168 46294
rect 254848 46170 254918 46226
rect 254974 46170 255042 46226
rect 255098 46170 255168 46226
rect 254848 46102 255168 46170
rect 254848 46046 254918 46102
rect 254974 46046 255042 46102
rect 255098 46046 255168 46102
rect 254848 45978 255168 46046
rect 254848 45922 254918 45978
rect 254974 45922 255042 45978
rect 255098 45922 255168 45978
rect 254848 45888 255168 45922
rect 285568 46350 285888 46384
rect 285568 46294 285638 46350
rect 285694 46294 285762 46350
rect 285818 46294 285888 46350
rect 285568 46226 285888 46294
rect 285568 46170 285638 46226
rect 285694 46170 285762 46226
rect 285818 46170 285888 46226
rect 285568 46102 285888 46170
rect 285568 46046 285638 46102
rect 285694 46046 285762 46102
rect 285818 46046 285888 46102
rect 285568 45978 285888 46046
rect 285568 45922 285638 45978
rect 285694 45922 285762 45978
rect 285818 45922 285888 45978
rect 285568 45888 285888 45922
rect 316288 46350 316608 46384
rect 316288 46294 316358 46350
rect 316414 46294 316482 46350
rect 316538 46294 316608 46350
rect 316288 46226 316608 46294
rect 316288 46170 316358 46226
rect 316414 46170 316482 46226
rect 316538 46170 316608 46226
rect 316288 46102 316608 46170
rect 316288 46046 316358 46102
rect 316414 46046 316482 46102
rect 316538 46046 316608 46102
rect 316288 45978 316608 46046
rect 316288 45922 316358 45978
rect 316414 45922 316482 45978
rect 316538 45922 316608 45978
rect 316288 45888 316608 45922
rect 347008 46350 347328 46384
rect 347008 46294 347078 46350
rect 347134 46294 347202 46350
rect 347258 46294 347328 46350
rect 347008 46226 347328 46294
rect 347008 46170 347078 46226
rect 347134 46170 347202 46226
rect 347258 46170 347328 46226
rect 347008 46102 347328 46170
rect 347008 46046 347078 46102
rect 347134 46046 347202 46102
rect 347258 46046 347328 46102
rect 347008 45978 347328 46046
rect 347008 45922 347078 45978
rect 347134 45922 347202 45978
rect 347258 45922 347328 45978
rect 347008 45888 347328 45922
rect 377728 46350 378048 46384
rect 377728 46294 377798 46350
rect 377854 46294 377922 46350
rect 377978 46294 378048 46350
rect 377728 46226 378048 46294
rect 377728 46170 377798 46226
rect 377854 46170 377922 46226
rect 377978 46170 378048 46226
rect 377728 46102 378048 46170
rect 377728 46046 377798 46102
rect 377854 46046 377922 46102
rect 377978 46046 378048 46102
rect 377728 45978 378048 46046
rect 377728 45922 377798 45978
rect 377854 45922 377922 45978
rect 377978 45922 378048 45978
rect 377728 45888 378048 45922
rect 408448 46350 408768 46384
rect 408448 46294 408518 46350
rect 408574 46294 408642 46350
rect 408698 46294 408768 46350
rect 408448 46226 408768 46294
rect 408448 46170 408518 46226
rect 408574 46170 408642 46226
rect 408698 46170 408768 46226
rect 408448 46102 408768 46170
rect 408448 46046 408518 46102
rect 408574 46046 408642 46102
rect 408698 46046 408768 46102
rect 408448 45978 408768 46046
rect 408448 45922 408518 45978
rect 408574 45922 408642 45978
rect 408698 45922 408768 45978
rect 408448 45888 408768 45922
rect 439168 46350 439488 46384
rect 439168 46294 439238 46350
rect 439294 46294 439362 46350
rect 439418 46294 439488 46350
rect 439168 46226 439488 46294
rect 439168 46170 439238 46226
rect 439294 46170 439362 46226
rect 439418 46170 439488 46226
rect 439168 46102 439488 46170
rect 439168 46046 439238 46102
rect 439294 46046 439362 46102
rect 439418 46046 439488 46102
rect 439168 45978 439488 46046
rect 439168 45922 439238 45978
rect 439294 45922 439362 45978
rect 439418 45922 439488 45978
rect 439168 45888 439488 45922
rect 469888 46350 470208 46384
rect 469888 46294 469958 46350
rect 470014 46294 470082 46350
rect 470138 46294 470208 46350
rect 469888 46226 470208 46294
rect 469888 46170 469958 46226
rect 470014 46170 470082 46226
rect 470138 46170 470208 46226
rect 469888 46102 470208 46170
rect 469888 46046 469958 46102
rect 470014 46046 470082 46102
rect 470138 46046 470208 46102
rect 469888 45978 470208 46046
rect 469888 45922 469958 45978
rect 470014 45922 470082 45978
rect 470138 45922 470208 45978
rect 469888 45888 470208 45922
rect 500608 46350 500928 46384
rect 500608 46294 500678 46350
rect 500734 46294 500802 46350
rect 500858 46294 500928 46350
rect 500608 46226 500928 46294
rect 500608 46170 500678 46226
rect 500734 46170 500802 46226
rect 500858 46170 500928 46226
rect 500608 46102 500928 46170
rect 500608 46046 500678 46102
rect 500734 46046 500802 46102
rect 500858 46046 500928 46102
rect 500608 45978 500928 46046
rect 500608 45922 500678 45978
rect 500734 45922 500802 45978
rect 500858 45922 500928 45978
rect 500608 45888 500928 45922
rect 24448 40350 24768 40384
rect 24448 40294 24518 40350
rect 24574 40294 24642 40350
rect 24698 40294 24768 40350
rect 24448 40226 24768 40294
rect 24448 40170 24518 40226
rect 24574 40170 24642 40226
rect 24698 40170 24768 40226
rect 24448 40102 24768 40170
rect 24448 40046 24518 40102
rect 24574 40046 24642 40102
rect 24698 40046 24768 40102
rect 24448 39978 24768 40046
rect 24448 39922 24518 39978
rect 24574 39922 24642 39978
rect 24698 39922 24768 39978
rect 24448 39888 24768 39922
rect 55168 40350 55488 40384
rect 55168 40294 55238 40350
rect 55294 40294 55362 40350
rect 55418 40294 55488 40350
rect 55168 40226 55488 40294
rect 55168 40170 55238 40226
rect 55294 40170 55362 40226
rect 55418 40170 55488 40226
rect 55168 40102 55488 40170
rect 55168 40046 55238 40102
rect 55294 40046 55362 40102
rect 55418 40046 55488 40102
rect 55168 39978 55488 40046
rect 55168 39922 55238 39978
rect 55294 39922 55362 39978
rect 55418 39922 55488 39978
rect 55168 39888 55488 39922
rect 85888 40350 86208 40384
rect 85888 40294 85958 40350
rect 86014 40294 86082 40350
rect 86138 40294 86208 40350
rect 85888 40226 86208 40294
rect 85888 40170 85958 40226
rect 86014 40170 86082 40226
rect 86138 40170 86208 40226
rect 85888 40102 86208 40170
rect 85888 40046 85958 40102
rect 86014 40046 86082 40102
rect 86138 40046 86208 40102
rect 85888 39978 86208 40046
rect 85888 39922 85958 39978
rect 86014 39922 86082 39978
rect 86138 39922 86208 39978
rect 85888 39888 86208 39922
rect 116608 40350 116928 40384
rect 116608 40294 116678 40350
rect 116734 40294 116802 40350
rect 116858 40294 116928 40350
rect 116608 40226 116928 40294
rect 116608 40170 116678 40226
rect 116734 40170 116802 40226
rect 116858 40170 116928 40226
rect 116608 40102 116928 40170
rect 116608 40046 116678 40102
rect 116734 40046 116802 40102
rect 116858 40046 116928 40102
rect 116608 39978 116928 40046
rect 116608 39922 116678 39978
rect 116734 39922 116802 39978
rect 116858 39922 116928 39978
rect 116608 39888 116928 39922
rect 147328 40350 147648 40384
rect 147328 40294 147398 40350
rect 147454 40294 147522 40350
rect 147578 40294 147648 40350
rect 147328 40226 147648 40294
rect 147328 40170 147398 40226
rect 147454 40170 147522 40226
rect 147578 40170 147648 40226
rect 147328 40102 147648 40170
rect 147328 40046 147398 40102
rect 147454 40046 147522 40102
rect 147578 40046 147648 40102
rect 147328 39978 147648 40046
rect 147328 39922 147398 39978
rect 147454 39922 147522 39978
rect 147578 39922 147648 39978
rect 147328 39888 147648 39922
rect 178048 40350 178368 40384
rect 178048 40294 178118 40350
rect 178174 40294 178242 40350
rect 178298 40294 178368 40350
rect 178048 40226 178368 40294
rect 178048 40170 178118 40226
rect 178174 40170 178242 40226
rect 178298 40170 178368 40226
rect 178048 40102 178368 40170
rect 178048 40046 178118 40102
rect 178174 40046 178242 40102
rect 178298 40046 178368 40102
rect 178048 39978 178368 40046
rect 178048 39922 178118 39978
rect 178174 39922 178242 39978
rect 178298 39922 178368 39978
rect 178048 39888 178368 39922
rect 208768 40350 209088 40384
rect 208768 40294 208838 40350
rect 208894 40294 208962 40350
rect 209018 40294 209088 40350
rect 208768 40226 209088 40294
rect 208768 40170 208838 40226
rect 208894 40170 208962 40226
rect 209018 40170 209088 40226
rect 208768 40102 209088 40170
rect 208768 40046 208838 40102
rect 208894 40046 208962 40102
rect 209018 40046 209088 40102
rect 208768 39978 209088 40046
rect 208768 39922 208838 39978
rect 208894 39922 208962 39978
rect 209018 39922 209088 39978
rect 208768 39888 209088 39922
rect 239488 40350 239808 40384
rect 239488 40294 239558 40350
rect 239614 40294 239682 40350
rect 239738 40294 239808 40350
rect 239488 40226 239808 40294
rect 239488 40170 239558 40226
rect 239614 40170 239682 40226
rect 239738 40170 239808 40226
rect 239488 40102 239808 40170
rect 239488 40046 239558 40102
rect 239614 40046 239682 40102
rect 239738 40046 239808 40102
rect 239488 39978 239808 40046
rect 239488 39922 239558 39978
rect 239614 39922 239682 39978
rect 239738 39922 239808 39978
rect 239488 39888 239808 39922
rect 270208 40350 270528 40384
rect 270208 40294 270278 40350
rect 270334 40294 270402 40350
rect 270458 40294 270528 40350
rect 270208 40226 270528 40294
rect 270208 40170 270278 40226
rect 270334 40170 270402 40226
rect 270458 40170 270528 40226
rect 270208 40102 270528 40170
rect 270208 40046 270278 40102
rect 270334 40046 270402 40102
rect 270458 40046 270528 40102
rect 270208 39978 270528 40046
rect 270208 39922 270278 39978
rect 270334 39922 270402 39978
rect 270458 39922 270528 39978
rect 270208 39888 270528 39922
rect 300928 40350 301248 40384
rect 300928 40294 300998 40350
rect 301054 40294 301122 40350
rect 301178 40294 301248 40350
rect 300928 40226 301248 40294
rect 300928 40170 300998 40226
rect 301054 40170 301122 40226
rect 301178 40170 301248 40226
rect 300928 40102 301248 40170
rect 300928 40046 300998 40102
rect 301054 40046 301122 40102
rect 301178 40046 301248 40102
rect 300928 39978 301248 40046
rect 300928 39922 300998 39978
rect 301054 39922 301122 39978
rect 301178 39922 301248 39978
rect 300928 39888 301248 39922
rect 331648 40350 331968 40384
rect 331648 40294 331718 40350
rect 331774 40294 331842 40350
rect 331898 40294 331968 40350
rect 331648 40226 331968 40294
rect 331648 40170 331718 40226
rect 331774 40170 331842 40226
rect 331898 40170 331968 40226
rect 331648 40102 331968 40170
rect 331648 40046 331718 40102
rect 331774 40046 331842 40102
rect 331898 40046 331968 40102
rect 331648 39978 331968 40046
rect 331648 39922 331718 39978
rect 331774 39922 331842 39978
rect 331898 39922 331968 39978
rect 331648 39888 331968 39922
rect 362368 40350 362688 40384
rect 362368 40294 362438 40350
rect 362494 40294 362562 40350
rect 362618 40294 362688 40350
rect 362368 40226 362688 40294
rect 362368 40170 362438 40226
rect 362494 40170 362562 40226
rect 362618 40170 362688 40226
rect 362368 40102 362688 40170
rect 362368 40046 362438 40102
rect 362494 40046 362562 40102
rect 362618 40046 362688 40102
rect 362368 39978 362688 40046
rect 362368 39922 362438 39978
rect 362494 39922 362562 39978
rect 362618 39922 362688 39978
rect 362368 39888 362688 39922
rect 393088 40350 393408 40384
rect 393088 40294 393158 40350
rect 393214 40294 393282 40350
rect 393338 40294 393408 40350
rect 393088 40226 393408 40294
rect 393088 40170 393158 40226
rect 393214 40170 393282 40226
rect 393338 40170 393408 40226
rect 393088 40102 393408 40170
rect 393088 40046 393158 40102
rect 393214 40046 393282 40102
rect 393338 40046 393408 40102
rect 393088 39978 393408 40046
rect 393088 39922 393158 39978
rect 393214 39922 393282 39978
rect 393338 39922 393408 39978
rect 393088 39888 393408 39922
rect 423808 40350 424128 40384
rect 423808 40294 423878 40350
rect 423934 40294 424002 40350
rect 424058 40294 424128 40350
rect 423808 40226 424128 40294
rect 423808 40170 423878 40226
rect 423934 40170 424002 40226
rect 424058 40170 424128 40226
rect 423808 40102 424128 40170
rect 423808 40046 423878 40102
rect 423934 40046 424002 40102
rect 424058 40046 424128 40102
rect 423808 39978 424128 40046
rect 423808 39922 423878 39978
rect 423934 39922 424002 39978
rect 424058 39922 424128 39978
rect 423808 39888 424128 39922
rect 454528 40350 454848 40384
rect 454528 40294 454598 40350
rect 454654 40294 454722 40350
rect 454778 40294 454848 40350
rect 454528 40226 454848 40294
rect 454528 40170 454598 40226
rect 454654 40170 454722 40226
rect 454778 40170 454848 40226
rect 454528 40102 454848 40170
rect 454528 40046 454598 40102
rect 454654 40046 454722 40102
rect 454778 40046 454848 40102
rect 454528 39978 454848 40046
rect 454528 39922 454598 39978
rect 454654 39922 454722 39978
rect 454778 39922 454848 39978
rect 454528 39888 454848 39922
rect 485248 40350 485568 40384
rect 485248 40294 485318 40350
rect 485374 40294 485442 40350
rect 485498 40294 485568 40350
rect 485248 40226 485568 40294
rect 485248 40170 485318 40226
rect 485374 40170 485442 40226
rect 485498 40170 485568 40226
rect 485248 40102 485568 40170
rect 485248 40046 485318 40102
rect 485374 40046 485442 40102
rect 485498 40046 485568 40102
rect 485248 39978 485568 40046
rect 485248 39922 485318 39978
rect 485374 39922 485442 39978
rect 485498 39922 485568 39978
rect 485248 39888 485568 39922
rect 515968 40350 516288 40384
rect 515968 40294 516038 40350
rect 516094 40294 516162 40350
rect 516218 40294 516288 40350
rect 515968 40226 516288 40294
rect 515968 40170 516038 40226
rect 516094 40170 516162 40226
rect 516218 40170 516288 40226
rect 515968 40102 516288 40170
rect 515968 40046 516038 40102
rect 516094 40046 516162 40102
rect 516218 40046 516288 40102
rect 515968 39978 516288 40046
rect 515968 39922 516038 39978
rect 516094 39922 516162 39978
rect 516218 39922 516288 39978
rect 515968 39888 516288 39922
rect 525154 40350 525774 57922
rect 525154 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 525774 40350
rect 525154 40226 525774 40294
rect 525154 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 525774 40226
rect 525154 40102 525774 40170
rect 525154 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 525774 40102
rect 525154 39978 525774 40046
rect 525154 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 525774 39978
rect 6874 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 7494 28350
rect 6874 28226 7494 28294
rect 6874 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 7494 28226
rect 6874 28102 7494 28170
rect 6874 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 7494 28102
rect 6874 27978 7494 28046
rect 6874 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 7494 27978
rect 6874 10350 7494 27922
rect 39808 28350 40128 28384
rect 39808 28294 39878 28350
rect 39934 28294 40002 28350
rect 40058 28294 40128 28350
rect 39808 28226 40128 28294
rect 39808 28170 39878 28226
rect 39934 28170 40002 28226
rect 40058 28170 40128 28226
rect 39808 28102 40128 28170
rect 39808 28046 39878 28102
rect 39934 28046 40002 28102
rect 40058 28046 40128 28102
rect 39808 27978 40128 28046
rect 39808 27922 39878 27978
rect 39934 27922 40002 27978
rect 40058 27922 40128 27978
rect 39808 27888 40128 27922
rect 70528 28350 70848 28384
rect 70528 28294 70598 28350
rect 70654 28294 70722 28350
rect 70778 28294 70848 28350
rect 70528 28226 70848 28294
rect 70528 28170 70598 28226
rect 70654 28170 70722 28226
rect 70778 28170 70848 28226
rect 70528 28102 70848 28170
rect 70528 28046 70598 28102
rect 70654 28046 70722 28102
rect 70778 28046 70848 28102
rect 70528 27978 70848 28046
rect 70528 27922 70598 27978
rect 70654 27922 70722 27978
rect 70778 27922 70848 27978
rect 70528 27888 70848 27922
rect 101248 28350 101568 28384
rect 101248 28294 101318 28350
rect 101374 28294 101442 28350
rect 101498 28294 101568 28350
rect 101248 28226 101568 28294
rect 101248 28170 101318 28226
rect 101374 28170 101442 28226
rect 101498 28170 101568 28226
rect 101248 28102 101568 28170
rect 101248 28046 101318 28102
rect 101374 28046 101442 28102
rect 101498 28046 101568 28102
rect 101248 27978 101568 28046
rect 101248 27922 101318 27978
rect 101374 27922 101442 27978
rect 101498 27922 101568 27978
rect 101248 27888 101568 27922
rect 131968 28350 132288 28384
rect 131968 28294 132038 28350
rect 132094 28294 132162 28350
rect 132218 28294 132288 28350
rect 131968 28226 132288 28294
rect 131968 28170 132038 28226
rect 132094 28170 132162 28226
rect 132218 28170 132288 28226
rect 131968 28102 132288 28170
rect 131968 28046 132038 28102
rect 132094 28046 132162 28102
rect 132218 28046 132288 28102
rect 131968 27978 132288 28046
rect 131968 27922 132038 27978
rect 132094 27922 132162 27978
rect 132218 27922 132288 27978
rect 131968 27888 132288 27922
rect 162688 28350 163008 28384
rect 162688 28294 162758 28350
rect 162814 28294 162882 28350
rect 162938 28294 163008 28350
rect 162688 28226 163008 28294
rect 162688 28170 162758 28226
rect 162814 28170 162882 28226
rect 162938 28170 163008 28226
rect 162688 28102 163008 28170
rect 162688 28046 162758 28102
rect 162814 28046 162882 28102
rect 162938 28046 163008 28102
rect 162688 27978 163008 28046
rect 162688 27922 162758 27978
rect 162814 27922 162882 27978
rect 162938 27922 163008 27978
rect 162688 27888 163008 27922
rect 193408 28350 193728 28384
rect 193408 28294 193478 28350
rect 193534 28294 193602 28350
rect 193658 28294 193728 28350
rect 193408 28226 193728 28294
rect 193408 28170 193478 28226
rect 193534 28170 193602 28226
rect 193658 28170 193728 28226
rect 193408 28102 193728 28170
rect 193408 28046 193478 28102
rect 193534 28046 193602 28102
rect 193658 28046 193728 28102
rect 193408 27978 193728 28046
rect 193408 27922 193478 27978
rect 193534 27922 193602 27978
rect 193658 27922 193728 27978
rect 193408 27888 193728 27922
rect 224128 28350 224448 28384
rect 224128 28294 224198 28350
rect 224254 28294 224322 28350
rect 224378 28294 224448 28350
rect 224128 28226 224448 28294
rect 224128 28170 224198 28226
rect 224254 28170 224322 28226
rect 224378 28170 224448 28226
rect 224128 28102 224448 28170
rect 224128 28046 224198 28102
rect 224254 28046 224322 28102
rect 224378 28046 224448 28102
rect 224128 27978 224448 28046
rect 224128 27922 224198 27978
rect 224254 27922 224322 27978
rect 224378 27922 224448 27978
rect 224128 27888 224448 27922
rect 254848 28350 255168 28384
rect 254848 28294 254918 28350
rect 254974 28294 255042 28350
rect 255098 28294 255168 28350
rect 254848 28226 255168 28294
rect 254848 28170 254918 28226
rect 254974 28170 255042 28226
rect 255098 28170 255168 28226
rect 254848 28102 255168 28170
rect 254848 28046 254918 28102
rect 254974 28046 255042 28102
rect 255098 28046 255168 28102
rect 254848 27978 255168 28046
rect 254848 27922 254918 27978
rect 254974 27922 255042 27978
rect 255098 27922 255168 27978
rect 254848 27888 255168 27922
rect 285568 28350 285888 28384
rect 285568 28294 285638 28350
rect 285694 28294 285762 28350
rect 285818 28294 285888 28350
rect 285568 28226 285888 28294
rect 285568 28170 285638 28226
rect 285694 28170 285762 28226
rect 285818 28170 285888 28226
rect 285568 28102 285888 28170
rect 285568 28046 285638 28102
rect 285694 28046 285762 28102
rect 285818 28046 285888 28102
rect 285568 27978 285888 28046
rect 285568 27922 285638 27978
rect 285694 27922 285762 27978
rect 285818 27922 285888 27978
rect 285568 27888 285888 27922
rect 316288 28350 316608 28384
rect 316288 28294 316358 28350
rect 316414 28294 316482 28350
rect 316538 28294 316608 28350
rect 316288 28226 316608 28294
rect 316288 28170 316358 28226
rect 316414 28170 316482 28226
rect 316538 28170 316608 28226
rect 316288 28102 316608 28170
rect 316288 28046 316358 28102
rect 316414 28046 316482 28102
rect 316538 28046 316608 28102
rect 316288 27978 316608 28046
rect 316288 27922 316358 27978
rect 316414 27922 316482 27978
rect 316538 27922 316608 27978
rect 316288 27888 316608 27922
rect 347008 28350 347328 28384
rect 347008 28294 347078 28350
rect 347134 28294 347202 28350
rect 347258 28294 347328 28350
rect 347008 28226 347328 28294
rect 347008 28170 347078 28226
rect 347134 28170 347202 28226
rect 347258 28170 347328 28226
rect 347008 28102 347328 28170
rect 347008 28046 347078 28102
rect 347134 28046 347202 28102
rect 347258 28046 347328 28102
rect 347008 27978 347328 28046
rect 347008 27922 347078 27978
rect 347134 27922 347202 27978
rect 347258 27922 347328 27978
rect 347008 27888 347328 27922
rect 377728 28350 378048 28384
rect 377728 28294 377798 28350
rect 377854 28294 377922 28350
rect 377978 28294 378048 28350
rect 377728 28226 378048 28294
rect 377728 28170 377798 28226
rect 377854 28170 377922 28226
rect 377978 28170 378048 28226
rect 377728 28102 378048 28170
rect 377728 28046 377798 28102
rect 377854 28046 377922 28102
rect 377978 28046 378048 28102
rect 377728 27978 378048 28046
rect 377728 27922 377798 27978
rect 377854 27922 377922 27978
rect 377978 27922 378048 27978
rect 377728 27888 378048 27922
rect 408448 28350 408768 28384
rect 408448 28294 408518 28350
rect 408574 28294 408642 28350
rect 408698 28294 408768 28350
rect 408448 28226 408768 28294
rect 408448 28170 408518 28226
rect 408574 28170 408642 28226
rect 408698 28170 408768 28226
rect 408448 28102 408768 28170
rect 408448 28046 408518 28102
rect 408574 28046 408642 28102
rect 408698 28046 408768 28102
rect 408448 27978 408768 28046
rect 408448 27922 408518 27978
rect 408574 27922 408642 27978
rect 408698 27922 408768 27978
rect 408448 27888 408768 27922
rect 439168 28350 439488 28384
rect 439168 28294 439238 28350
rect 439294 28294 439362 28350
rect 439418 28294 439488 28350
rect 439168 28226 439488 28294
rect 439168 28170 439238 28226
rect 439294 28170 439362 28226
rect 439418 28170 439488 28226
rect 439168 28102 439488 28170
rect 439168 28046 439238 28102
rect 439294 28046 439362 28102
rect 439418 28046 439488 28102
rect 439168 27978 439488 28046
rect 439168 27922 439238 27978
rect 439294 27922 439362 27978
rect 439418 27922 439488 27978
rect 439168 27888 439488 27922
rect 469888 28350 470208 28384
rect 469888 28294 469958 28350
rect 470014 28294 470082 28350
rect 470138 28294 470208 28350
rect 469888 28226 470208 28294
rect 469888 28170 469958 28226
rect 470014 28170 470082 28226
rect 470138 28170 470208 28226
rect 469888 28102 470208 28170
rect 469888 28046 469958 28102
rect 470014 28046 470082 28102
rect 470138 28046 470208 28102
rect 469888 27978 470208 28046
rect 469888 27922 469958 27978
rect 470014 27922 470082 27978
rect 470138 27922 470208 27978
rect 469888 27888 470208 27922
rect 500608 28350 500928 28384
rect 500608 28294 500678 28350
rect 500734 28294 500802 28350
rect 500858 28294 500928 28350
rect 500608 28226 500928 28294
rect 500608 28170 500678 28226
rect 500734 28170 500802 28226
rect 500858 28170 500928 28226
rect 500608 28102 500928 28170
rect 500608 28046 500678 28102
rect 500734 28046 500802 28102
rect 500858 28046 500928 28102
rect 500608 27978 500928 28046
rect 500608 27922 500678 27978
rect 500734 27922 500802 27978
rect 500858 27922 500928 27978
rect 500608 27888 500928 27922
rect 525154 22350 525774 39922
rect 525154 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 525774 22350
rect 525154 22226 525774 22294
rect 525154 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 525774 22226
rect 525154 22102 525774 22170
rect 525154 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 525774 22102
rect 525154 21978 525774 22046
rect 525154 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 525774 21978
rect 6874 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 7494 10350
rect 6874 10226 7494 10294
rect 6874 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 7494 10226
rect 6874 10102 7494 10170
rect 6874 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 7494 10102
rect 6874 9978 7494 10046
rect 6874 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 7494 9978
rect 6874 -1120 7494 9922
rect 6874 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 7494 -1120
rect 6874 -1244 7494 -1176
rect 6874 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 7494 -1244
rect 6874 -1368 7494 -1300
rect 6874 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 7494 -1368
rect 6874 -1492 7494 -1424
rect 6874 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 7494 -1492
rect 6874 -1644 7494 -1548
rect 21154 4350 21774 18186
rect 21154 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 21774 4350
rect 21154 4226 21774 4294
rect 21154 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 21774 4226
rect 21154 4102 21774 4170
rect 21154 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 21774 4102
rect 21154 3978 21774 4046
rect 21154 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 21774 3978
rect 21154 -160 21774 3922
rect 21154 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 21774 -160
rect 21154 -284 21774 -216
rect 21154 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 21774 -284
rect 21154 -408 21774 -340
rect 21154 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 21774 -408
rect 21154 -532 21774 -464
rect 21154 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 21774 -532
rect 21154 -1644 21774 -588
rect 24874 10350 25494 18186
rect 24874 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 25494 10350
rect 24874 10226 25494 10294
rect 24874 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 25494 10226
rect 24874 10102 25494 10170
rect 24874 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 25494 10102
rect 24874 9978 25494 10046
rect 24874 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 25494 9978
rect 24874 -1120 25494 9922
rect 24874 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 25494 -1120
rect 24874 -1244 25494 -1176
rect 24874 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 25494 -1244
rect 24874 -1368 25494 -1300
rect 24874 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 25494 -1368
rect 24874 -1492 25494 -1424
rect 24874 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 25494 -1492
rect 24874 -1644 25494 -1548
rect 39154 4350 39774 18186
rect 39154 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 39774 4350
rect 39154 4226 39774 4294
rect 39154 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 39774 4226
rect 39154 4102 39774 4170
rect 39154 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 39774 4102
rect 39154 3978 39774 4046
rect 39154 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 39774 3978
rect 39154 -160 39774 3922
rect 39154 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 39774 -160
rect 39154 -284 39774 -216
rect 39154 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 39774 -284
rect 39154 -408 39774 -340
rect 39154 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 39774 -408
rect 39154 -532 39774 -464
rect 39154 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 39774 -532
rect 39154 -1644 39774 -588
rect 42874 10350 43494 18186
rect 42874 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 43494 10350
rect 42874 10226 43494 10294
rect 42874 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 43494 10226
rect 42874 10102 43494 10170
rect 42874 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 43494 10102
rect 42874 9978 43494 10046
rect 42874 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 43494 9978
rect 42874 -1120 43494 9922
rect 42874 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 43494 -1120
rect 42874 -1244 43494 -1176
rect 42874 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 43494 -1244
rect 42874 -1368 43494 -1300
rect 42874 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 43494 -1368
rect 42874 -1492 43494 -1424
rect 42874 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 43494 -1492
rect 42874 -1644 43494 -1548
rect 57154 4350 57774 18186
rect 57154 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 57774 4350
rect 57154 4226 57774 4294
rect 57154 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 57774 4226
rect 57154 4102 57774 4170
rect 57154 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 57774 4102
rect 57154 3978 57774 4046
rect 57154 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 57774 3978
rect 57154 -160 57774 3922
rect 57154 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 57774 -160
rect 57154 -284 57774 -216
rect 57154 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 57774 -284
rect 57154 -408 57774 -340
rect 57154 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 57774 -408
rect 57154 -532 57774 -464
rect 57154 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 57774 -532
rect 57154 -1644 57774 -588
rect 60874 10350 61494 18186
rect 60874 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 61494 10350
rect 60874 10226 61494 10294
rect 60874 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 61494 10226
rect 60874 10102 61494 10170
rect 60874 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 61494 10102
rect 60874 9978 61494 10046
rect 60874 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 61494 9978
rect 60874 -1120 61494 9922
rect 60874 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 61494 -1120
rect 60874 -1244 61494 -1176
rect 60874 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 61494 -1244
rect 60874 -1368 61494 -1300
rect 60874 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 61494 -1368
rect 60874 -1492 61494 -1424
rect 60874 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 61494 -1492
rect 60874 -1644 61494 -1548
rect 75154 4350 75774 18186
rect 75154 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 75774 4350
rect 75154 4226 75774 4294
rect 75154 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 75774 4226
rect 75154 4102 75774 4170
rect 75154 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 75774 4102
rect 75154 3978 75774 4046
rect 75154 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 75774 3978
rect 75154 -160 75774 3922
rect 75154 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 75774 -160
rect 75154 -284 75774 -216
rect 75154 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 75774 -284
rect 75154 -408 75774 -340
rect 75154 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 75774 -408
rect 75154 -532 75774 -464
rect 75154 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 75774 -532
rect 75154 -1644 75774 -588
rect 78874 10350 79494 18186
rect 78874 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 79494 10350
rect 78874 10226 79494 10294
rect 78874 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 79494 10226
rect 78874 10102 79494 10170
rect 78874 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 79494 10102
rect 78874 9978 79494 10046
rect 78874 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 79494 9978
rect 78874 -1120 79494 9922
rect 78874 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 79494 -1120
rect 78874 -1244 79494 -1176
rect 78874 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 79494 -1244
rect 78874 -1368 79494 -1300
rect 78874 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 79494 -1368
rect 78874 -1492 79494 -1424
rect 78874 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 79494 -1492
rect 78874 -1644 79494 -1548
rect 93154 4350 93774 18186
rect 93154 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 93774 4350
rect 93154 4226 93774 4294
rect 93154 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 93774 4226
rect 93154 4102 93774 4170
rect 93154 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 93774 4102
rect 93154 3978 93774 4046
rect 93154 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 93774 3978
rect 93154 -160 93774 3922
rect 93154 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 93774 -160
rect 93154 -284 93774 -216
rect 93154 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 93774 -284
rect 93154 -408 93774 -340
rect 93154 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 93774 -408
rect 93154 -532 93774 -464
rect 93154 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 93774 -532
rect 93154 -1644 93774 -588
rect 96874 10350 97494 18186
rect 96874 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 97494 10350
rect 96874 10226 97494 10294
rect 96874 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 97494 10226
rect 96874 10102 97494 10170
rect 96874 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 97494 10102
rect 96874 9978 97494 10046
rect 96874 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 97494 9978
rect 96874 -1120 97494 9922
rect 96874 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 97494 -1120
rect 96874 -1244 97494 -1176
rect 96874 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 97494 -1244
rect 96874 -1368 97494 -1300
rect 96874 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 97494 -1368
rect 96874 -1492 97494 -1424
rect 96874 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 97494 -1492
rect 96874 -1644 97494 -1548
rect 111154 4350 111774 18186
rect 111154 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 111774 4350
rect 111154 4226 111774 4294
rect 111154 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 111774 4226
rect 111154 4102 111774 4170
rect 111154 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 111774 4102
rect 111154 3978 111774 4046
rect 111154 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 111774 3978
rect 111154 -160 111774 3922
rect 111154 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 111774 -160
rect 111154 -284 111774 -216
rect 111154 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 111774 -284
rect 111154 -408 111774 -340
rect 111154 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 111774 -408
rect 111154 -532 111774 -464
rect 111154 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 111774 -532
rect 111154 -1644 111774 -588
rect 114874 10350 115494 18186
rect 114874 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 115494 10350
rect 114874 10226 115494 10294
rect 114874 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 115494 10226
rect 114874 10102 115494 10170
rect 114874 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 115494 10102
rect 114874 9978 115494 10046
rect 114874 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 115494 9978
rect 114874 -1120 115494 9922
rect 114874 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 115494 -1120
rect 114874 -1244 115494 -1176
rect 114874 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 115494 -1244
rect 114874 -1368 115494 -1300
rect 114874 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 115494 -1368
rect 114874 -1492 115494 -1424
rect 114874 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 115494 -1492
rect 114874 -1644 115494 -1548
rect 129154 4350 129774 18186
rect 129154 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 129774 4350
rect 129154 4226 129774 4294
rect 129154 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 129774 4226
rect 129154 4102 129774 4170
rect 129154 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 129774 4102
rect 129154 3978 129774 4046
rect 129154 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 129774 3978
rect 129154 -160 129774 3922
rect 129154 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 129774 -160
rect 129154 -284 129774 -216
rect 129154 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 129774 -284
rect 129154 -408 129774 -340
rect 129154 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 129774 -408
rect 129154 -532 129774 -464
rect 129154 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 129774 -532
rect 129154 -1644 129774 -588
rect 132874 10350 133494 18186
rect 132874 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 133494 10350
rect 132874 10226 133494 10294
rect 132874 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 133494 10226
rect 132874 10102 133494 10170
rect 132874 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 133494 10102
rect 132874 9978 133494 10046
rect 132874 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 133494 9978
rect 132874 -1120 133494 9922
rect 132874 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 133494 -1120
rect 132874 -1244 133494 -1176
rect 132874 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 133494 -1244
rect 132874 -1368 133494 -1300
rect 132874 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 133494 -1368
rect 132874 -1492 133494 -1424
rect 132874 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 133494 -1492
rect 132874 -1644 133494 -1548
rect 147154 4350 147774 18186
rect 147154 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 147774 4350
rect 147154 4226 147774 4294
rect 147154 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 147774 4226
rect 147154 4102 147774 4170
rect 147154 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 147774 4102
rect 147154 3978 147774 4046
rect 147154 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 147774 3978
rect 147154 -160 147774 3922
rect 147154 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 147774 -160
rect 147154 -284 147774 -216
rect 147154 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 147774 -284
rect 147154 -408 147774 -340
rect 147154 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 147774 -408
rect 147154 -532 147774 -464
rect 147154 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 147774 -532
rect 147154 -1644 147774 -588
rect 150874 10350 151494 18186
rect 150874 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 151494 10350
rect 150874 10226 151494 10294
rect 150874 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 151494 10226
rect 150874 10102 151494 10170
rect 150874 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 151494 10102
rect 150874 9978 151494 10046
rect 150874 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 151494 9978
rect 150874 -1120 151494 9922
rect 150874 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 151494 -1120
rect 150874 -1244 151494 -1176
rect 150874 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 151494 -1244
rect 150874 -1368 151494 -1300
rect 150874 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 151494 -1368
rect 150874 -1492 151494 -1424
rect 150874 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 151494 -1492
rect 150874 -1644 151494 -1548
rect 165154 4350 165774 18186
rect 165154 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 165774 4350
rect 165154 4226 165774 4294
rect 165154 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 165774 4226
rect 165154 4102 165774 4170
rect 165154 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 165774 4102
rect 165154 3978 165774 4046
rect 165154 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 165774 3978
rect 165154 -160 165774 3922
rect 165154 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 165774 -160
rect 165154 -284 165774 -216
rect 165154 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 165774 -284
rect 165154 -408 165774 -340
rect 165154 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 165774 -408
rect 165154 -532 165774 -464
rect 165154 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 165774 -532
rect 165154 -1644 165774 -588
rect 168874 10350 169494 18186
rect 168874 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 169494 10350
rect 168874 10226 169494 10294
rect 168874 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 169494 10226
rect 168874 10102 169494 10170
rect 168874 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 169494 10102
rect 168874 9978 169494 10046
rect 168874 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 169494 9978
rect 168874 -1120 169494 9922
rect 168874 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 169494 -1120
rect 168874 -1244 169494 -1176
rect 168874 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 169494 -1244
rect 168874 -1368 169494 -1300
rect 168874 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 169494 -1368
rect 168874 -1492 169494 -1424
rect 168874 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 169494 -1492
rect 168874 -1644 169494 -1548
rect 183154 4350 183774 18186
rect 183154 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 183774 4350
rect 183154 4226 183774 4294
rect 183154 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 183774 4226
rect 183154 4102 183774 4170
rect 183154 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 183774 4102
rect 183154 3978 183774 4046
rect 183154 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 183774 3978
rect 183154 -160 183774 3922
rect 183154 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 183774 -160
rect 183154 -284 183774 -216
rect 183154 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 183774 -284
rect 183154 -408 183774 -340
rect 183154 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 183774 -408
rect 183154 -532 183774 -464
rect 183154 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 183774 -532
rect 183154 -1644 183774 -588
rect 186874 10350 187494 18186
rect 186874 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 187494 10350
rect 186874 10226 187494 10294
rect 186874 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 187494 10226
rect 186874 10102 187494 10170
rect 186874 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 187494 10102
rect 186874 9978 187494 10046
rect 186874 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 187494 9978
rect 186874 -1120 187494 9922
rect 186874 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 187494 -1120
rect 186874 -1244 187494 -1176
rect 186874 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 187494 -1244
rect 186874 -1368 187494 -1300
rect 186874 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 187494 -1368
rect 186874 -1492 187494 -1424
rect 186874 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 187494 -1492
rect 186874 -1644 187494 -1548
rect 201154 4350 201774 18186
rect 201154 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 201774 4350
rect 201154 4226 201774 4294
rect 201154 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 201774 4226
rect 201154 4102 201774 4170
rect 201154 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 201774 4102
rect 201154 3978 201774 4046
rect 201154 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 201774 3978
rect 201154 -160 201774 3922
rect 201154 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 201774 -160
rect 201154 -284 201774 -216
rect 201154 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 201774 -284
rect 201154 -408 201774 -340
rect 201154 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 201774 -408
rect 201154 -532 201774 -464
rect 201154 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 201774 -532
rect 201154 -1644 201774 -588
rect 204874 10350 205494 18186
rect 204874 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 205494 10350
rect 204874 10226 205494 10294
rect 204874 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 205494 10226
rect 204874 10102 205494 10170
rect 204874 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 205494 10102
rect 204874 9978 205494 10046
rect 204874 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 205494 9978
rect 204874 -1120 205494 9922
rect 204874 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 205494 -1120
rect 204874 -1244 205494 -1176
rect 204874 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 205494 -1244
rect 204874 -1368 205494 -1300
rect 204874 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 205494 -1368
rect 204874 -1492 205494 -1424
rect 204874 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 205494 -1492
rect 204874 -1644 205494 -1548
rect 219154 4350 219774 18186
rect 219154 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 219774 4350
rect 219154 4226 219774 4294
rect 219154 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 219774 4226
rect 219154 4102 219774 4170
rect 219154 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 219774 4102
rect 219154 3978 219774 4046
rect 219154 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 219774 3978
rect 219154 -160 219774 3922
rect 219154 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 219774 -160
rect 219154 -284 219774 -216
rect 219154 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 219774 -284
rect 219154 -408 219774 -340
rect 219154 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 219774 -408
rect 219154 -532 219774 -464
rect 219154 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 219774 -532
rect 219154 -1644 219774 -588
rect 222874 10350 223494 18186
rect 222874 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 223494 10350
rect 222874 10226 223494 10294
rect 222874 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 223494 10226
rect 222874 10102 223494 10170
rect 222874 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 223494 10102
rect 222874 9978 223494 10046
rect 222874 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 223494 9978
rect 222874 -1120 223494 9922
rect 222874 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 223494 -1120
rect 222874 -1244 223494 -1176
rect 222874 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 223494 -1244
rect 222874 -1368 223494 -1300
rect 222874 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 223494 -1368
rect 222874 -1492 223494 -1424
rect 222874 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 223494 -1492
rect 222874 -1644 223494 -1548
rect 237154 4350 237774 18186
rect 237154 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 237774 4350
rect 237154 4226 237774 4294
rect 237154 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 237774 4226
rect 237154 4102 237774 4170
rect 237154 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 237774 4102
rect 237154 3978 237774 4046
rect 237154 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 237774 3978
rect 237154 -160 237774 3922
rect 237154 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 237774 -160
rect 237154 -284 237774 -216
rect 237154 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 237774 -284
rect 237154 -408 237774 -340
rect 237154 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 237774 -408
rect 237154 -532 237774 -464
rect 237154 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 237774 -532
rect 237154 -1644 237774 -588
rect 240874 10350 241494 18186
rect 240874 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 241494 10350
rect 240874 10226 241494 10294
rect 240874 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 241494 10226
rect 240874 10102 241494 10170
rect 240874 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 241494 10102
rect 240874 9978 241494 10046
rect 240874 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 241494 9978
rect 240874 -1120 241494 9922
rect 240874 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 241494 -1120
rect 240874 -1244 241494 -1176
rect 240874 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 241494 -1244
rect 240874 -1368 241494 -1300
rect 240874 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 241494 -1368
rect 240874 -1492 241494 -1424
rect 240874 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 241494 -1492
rect 240874 -1644 241494 -1548
rect 255154 4350 255774 18186
rect 255154 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 255774 4350
rect 255154 4226 255774 4294
rect 255154 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 255774 4226
rect 255154 4102 255774 4170
rect 255154 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 255774 4102
rect 255154 3978 255774 4046
rect 255154 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 255774 3978
rect 255154 -160 255774 3922
rect 255154 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 255774 -160
rect 255154 -284 255774 -216
rect 255154 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 255774 -284
rect 255154 -408 255774 -340
rect 255154 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 255774 -408
rect 255154 -532 255774 -464
rect 255154 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 255774 -532
rect 255154 -1644 255774 -588
rect 258874 10350 259494 18186
rect 258874 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 259494 10350
rect 258874 10226 259494 10294
rect 258874 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 259494 10226
rect 258874 10102 259494 10170
rect 258874 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 259494 10102
rect 258874 9978 259494 10046
rect 258874 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 259494 9978
rect 258874 -1120 259494 9922
rect 258874 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 259494 -1120
rect 258874 -1244 259494 -1176
rect 258874 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 259494 -1244
rect 258874 -1368 259494 -1300
rect 258874 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 259494 -1368
rect 258874 -1492 259494 -1424
rect 258874 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 259494 -1492
rect 258874 -1644 259494 -1548
rect 273154 4350 273774 18186
rect 273154 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 273774 4350
rect 273154 4226 273774 4294
rect 273154 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 273774 4226
rect 273154 4102 273774 4170
rect 273154 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 273774 4102
rect 273154 3978 273774 4046
rect 273154 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 273774 3978
rect 273154 -160 273774 3922
rect 273154 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 273774 -160
rect 273154 -284 273774 -216
rect 273154 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 273774 -284
rect 273154 -408 273774 -340
rect 273154 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 273774 -408
rect 273154 -532 273774 -464
rect 273154 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 273774 -532
rect 273154 -1644 273774 -588
rect 276874 10350 277494 18186
rect 276874 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 277494 10350
rect 276874 10226 277494 10294
rect 276874 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 277494 10226
rect 276874 10102 277494 10170
rect 276874 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 277494 10102
rect 276874 9978 277494 10046
rect 276874 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 277494 9978
rect 276874 -1120 277494 9922
rect 276874 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 277494 -1120
rect 276874 -1244 277494 -1176
rect 276874 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 277494 -1244
rect 276874 -1368 277494 -1300
rect 276874 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 277494 -1368
rect 276874 -1492 277494 -1424
rect 276874 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 277494 -1492
rect 276874 -1644 277494 -1548
rect 291154 4350 291774 18186
rect 291154 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 291774 4350
rect 291154 4226 291774 4294
rect 291154 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 291774 4226
rect 291154 4102 291774 4170
rect 291154 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 291774 4102
rect 291154 3978 291774 4046
rect 291154 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 291774 3978
rect 291154 -160 291774 3922
rect 291154 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 291774 -160
rect 291154 -284 291774 -216
rect 291154 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 291774 -284
rect 291154 -408 291774 -340
rect 291154 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 291774 -408
rect 291154 -532 291774 -464
rect 291154 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 291774 -532
rect 291154 -1644 291774 -588
rect 294874 10350 295494 18186
rect 294874 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 295494 10350
rect 294874 10226 295494 10294
rect 294874 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 295494 10226
rect 294874 10102 295494 10170
rect 294874 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 295494 10102
rect 294874 9978 295494 10046
rect 294874 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 295494 9978
rect 294874 -1120 295494 9922
rect 294874 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 295494 -1120
rect 294874 -1244 295494 -1176
rect 294874 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 295494 -1244
rect 294874 -1368 295494 -1300
rect 294874 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 295494 -1368
rect 294874 -1492 295494 -1424
rect 294874 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 295494 -1492
rect 294874 -1644 295494 -1548
rect 309154 4350 309774 18186
rect 309154 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 309774 4350
rect 309154 4226 309774 4294
rect 309154 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 309774 4226
rect 309154 4102 309774 4170
rect 309154 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 309774 4102
rect 309154 3978 309774 4046
rect 309154 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 309774 3978
rect 309154 -160 309774 3922
rect 309154 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 309774 -160
rect 309154 -284 309774 -216
rect 309154 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 309774 -284
rect 309154 -408 309774 -340
rect 309154 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 309774 -408
rect 309154 -532 309774 -464
rect 309154 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 309774 -532
rect 309154 -1644 309774 -588
rect 312874 10350 313494 18186
rect 312874 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 313494 10350
rect 312874 10226 313494 10294
rect 312874 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 313494 10226
rect 312874 10102 313494 10170
rect 312874 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 313494 10102
rect 312874 9978 313494 10046
rect 312874 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 313494 9978
rect 312874 -1120 313494 9922
rect 312874 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 313494 -1120
rect 312874 -1244 313494 -1176
rect 312874 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 313494 -1244
rect 312874 -1368 313494 -1300
rect 312874 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 313494 -1368
rect 312874 -1492 313494 -1424
rect 312874 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 313494 -1492
rect 312874 -1644 313494 -1548
rect 327154 4350 327774 18186
rect 327154 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 327774 4350
rect 327154 4226 327774 4294
rect 327154 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 327774 4226
rect 327154 4102 327774 4170
rect 327154 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 327774 4102
rect 327154 3978 327774 4046
rect 327154 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 327774 3978
rect 327154 -160 327774 3922
rect 327154 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 327774 -160
rect 327154 -284 327774 -216
rect 327154 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 327774 -284
rect 327154 -408 327774 -340
rect 327154 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 327774 -408
rect 327154 -532 327774 -464
rect 327154 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 327774 -532
rect 327154 -1644 327774 -588
rect 330874 10350 331494 18186
rect 330874 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 331494 10350
rect 330874 10226 331494 10294
rect 330874 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 331494 10226
rect 330874 10102 331494 10170
rect 330874 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 331494 10102
rect 330874 9978 331494 10046
rect 330874 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 331494 9978
rect 330874 -1120 331494 9922
rect 330874 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 331494 -1120
rect 330874 -1244 331494 -1176
rect 330874 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 331494 -1244
rect 330874 -1368 331494 -1300
rect 330874 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 331494 -1368
rect 330874 -1492 331494 -1424
rect 330874 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 331494 -1492
rect 330874 -1644 331494 -1548
rect 345154 4350 345774 18186
rect 345154 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 345774 4350
rect 345154 4226 345774 4294
rect 345154 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 345774 4226
rect 345154 4102 345774 4170
rect 345154 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 345774 4102
rect 345154 3978 345774 4046
rect 345154 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 345774 3978
rect 345154 -160 345774 3922
rect 345154 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 345774 -160
rect 345154 -284 345774 -216
rect 345154 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 345774 -284
rect 345154 -408 345774 -340
rect 345154 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 345774 -408
rect 345154 -532 345774 -464
rect 345154 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 345774 -532
rect 345154 -1644 345774 -588
rect 348874 10350 349494 18186
rect 348874 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 349494 10350
rect 348874 10226 349494 10294
rect 348874 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 349494 10226
rect 348874 10102 349494 10170
rect 348874 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 349494 10102
rect 348874 9978 349494 10046
rect 348874 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 349494 9978
rect 348874 -1120 349494 9922
rect 348874 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 349494 -1120
rect 348874 -1244 349494 -1176
rect 348874 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 349494 -1244
rect 348874 -1368 349494 -1300
rect 348874 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 349494 -1368
rect 348874 -1492 349494 -1424
rect 348874 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 349494 -1492
rect 348874 -1644 349494 -1548
rect 363154 4350 363774 18186
rect 363154 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 363774 4350
rect 363154 4226 363774 4294
rect 363154 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 363774 4226
rect 363154 4102 363774 4170
rect 363154 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 363774 4102
rect 363154 3978 363774 4046
rect 363154 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 363774 3978
rect 363154 -160 363774 3922
rect 363154 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 363774 -160
rect 363154 -284 363774 -216
rect 363154 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 363774 -284
rect 363154 -408 363774 -340
rect 363154 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 363774 -408
rect 363154 -532 363774 -464
rect 363154 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 363774 -532
rect 363154 -1644 363774 -588
rect 366874 10350 367494 18186
rect 366874 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 367494 10350
rect 366874 10226 367494 10294
rect 366874 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 367494 10226
rect 366874 10102 367494 10170
rect 366874 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 367494 10102
rect 366874 9978 367494 10046
rect 366874 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 367494 9978
rect 366874 -1120 367494 9922
rect 366874 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 367494 -1120
rect 366874 -1244 367494 -1176
rect 366874 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 367494 -1244
rect 366874 -1368 367494 -1300
rect 366874 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 367494 -1368
rect 366874 -1492 367494 -1424
rect 366874 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 367494 -1492
rect 366874 -1644 367494 -1548
rect 381154 4350 381774 18186
rect 381154 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 381774 4350
rect 381154 4226 381774 4294
rect 381154 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 381774 4226
rect 381154 4102 381774 4170
rect 381154 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 381774 4102
rect 381154 3978 381774 4046
rect 381154 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 381774 3978
rect 381154 -160 381774 3922
rect 381154 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 381774 -160
rect 381154 -284 381774 -216
rect 381154 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 381774 -284
rect 381154 -408 381774 -340
rect 381154 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 381774 -408
rect 381154 -532 381774 -464
rect 381154 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 381774 -532
rect 381154 -1644 381774 -588
rect 384874 10350 385494 18186
rect 384874 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 385494 10350
rect 384874 10226 385494 10294
rect 384874 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 385494 10226
rect 384874 10102 385494 10170
rect 384874 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 385494 10102
rect 384874 9978 385494 10046
rect 384874 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 385494 9978
rect 384874 -1120 385494 9922
rect 384874 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 385494 -1120
rect 384874 -1244 385494 -1176
rect 384874 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 385494 -1244
rect 384874 -1368 385494 -1300
rect 384874 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 385494 -1368
rect 384874 -1492 385494 -1424
rect 384874 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 385494 -1492
rect 384874 -1644 385494 -1548
rect 399154 4350 399774 18186
rect 399154 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 399774 4350
rect 399154 4226 399774 4294
rect 399154 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 399774 4226
rect 399154 4102 399774 4170
rect 399154 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 399774 4102
rect 399154 3978 399774 4046
rect 399154 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 399774 3978
rect 399154 -160 399774 3922
rect 399154 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 399774 -160
rect 399154 -284 399774 -216
rect 399154 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 399774 -284
rect 399154 -408 399774 -340
rect 399154 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 399774 -408
rect 399154 -532 399774 -464
rect 399154 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 399774 -532
rect 399154 -1644 399774 -588
rect 402874 10350 403494 18186
rect 402874 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 403494 10350
rect 402874 10226 403494 10294
rect 402874 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 403494 10226
rect 402874 10102 403494 10170
rect 402874 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 403494 10102
rect 402874 9978 403494 10046
rect 402874 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 403494 9978
rect 402874 -1120 403494 9922
rect 402874 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 403494 -1120
rect 402874 -1244 403494 -1176
rect 402874 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 403494 -1244
rect 402874 -1368 403494 -1300
rect 402874 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 403494 -1368
rect 402874 -1492 403494 -1424
rect 402874 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 403494 -1492
rect 402874 -1644 403494 -1548
rect 417154 4350 417774 18186
rect 417154 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 417774 4350
rect 417154 4226 417774 4294
rect 417154 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 417774 4226
rect 417154 4102 417774 4170
rect 417154 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 417774 4102
rect 417154 3978 417774 4046
rect 417154 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 417774 3978
rect 417154 -160 417774 3922
rect 417154 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 417774 -160
rect 417154 -284 417774 -216
rect 417154 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 417774 -284
rect 417154 -408 417774 -340
rect 417154 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 417774 -408
rect 417154 -532 417774 -464
rect 417154 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 417774 -532
rect 417154 -1644 417774 -588
rect 420874 10350 421494 18186
rect 420874 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 421494 10350
rect 420874 10226 421494 10294
rect 420874 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 421494 10226
rect 420874 10102 421494 10170
rect 420874 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 421494 10102
rect 420874 9978 421494 10046
rect 420874 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 421494 9978
rect 420874 -1120 421494 9922
rect 420874 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 421494 -1120
rect 420874 -1244 421494 -1176
rect 420874 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 421494 -1244
rect 420874 -1368 421494 -1300
rect 420874 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 421494 -1368
rect 420874 -1492 421494 -1424
rect 420874 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 421494 -1492
rect 420874 -1644 421494 -1548
rect 435154 4350 435774 18186
rect 435154 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 435774 4350
rect 435154 4226 435774 4294
rect 435154 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 435774 4226
rect 435154 4102 435774 4170
rect 435154 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 435774 4102
rect 435154 3978 435774 4046
rect 435154 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 435774 3978
rect 435154 -160 435774 3922
rect 435154 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 435774 -160
rect 435154 -284 435774 -216
rect 435154 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 435774 -284
rect 435154 -408 435774 -340
rect 435154 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 435774 -408
rect 435154 -532 435774 -464
rect 435154 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 435774 -532
rect 435154 -1644 435774 -588
rect 438874 10350 439494 18186
rect 438874 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 439494 10350
rect 438874 10226 439494 10294
rect 438874 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 439494 10226
rect 438874 10102 439494 10170
rect 438874 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 439494 10102
rect 438874 9978 439494 10046
rect 438874 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 439494 9978
rect 438874 -1120 439494 9922
rect 438874 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 439494 -1120
rect 438874 -1244 439494 -1176
rect 438874 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 439494 -1244
rect 438874 -1368 439494 -1300
rect 438874 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 439494 -1368
rect 438874 -1492 439494 -1424
rect 438874 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 439494 -1492
rect 438874 -1644 439494 -1548
rect 453154 4350 453774 18186
rect 453154 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 453774 4350
rect 453154 4226 453774 4294
rect 453154 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 453774 4226
rect 453154 4102 453774 4170
rect 453154 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 453774 4102
rect 453154 3978 453774 4046
rect 453154 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 453774 3978
rect 453154 -160 453774 3922
rect 453154 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 453774 -160
rect 453154 -284 453774 -216
rect 453154 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 453774 -284
rect 453154 -408 453774 -340
rect 453154 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 453774 -408
rect 453154 -532 453774 -464
rect 453154 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 453774 -532
rect 453154 -1644 453774 -588
rect 456874 10350 457494 18186
rect 456874 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 457494 10350
rect 456874 10226 457494 10294
rect 456874 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 457494 10226
rect 456874 10102 457494 10170
rect 456874 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 457494 10102
rect 456874 9978 457494 10046
rect 456874 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 457494 9978
rect 456874 -1120 457494 9922
rect 456874 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 457494 -1120
rect 456874 -1244 457494 -1176
rect 456874 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 457494 -1244
rect 456874 -1368 457494 -1300
rect 456874 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 457494 -1368
rect 456874 -1492 457494 -1424
rect 456874 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 457494 -1492
rect 456874 -1644 457494 -1548
rect 471154 4350 471774 18186
rect 471154 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 471774 4350
rect 471154 4226 471774 4294
rect 471154 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 471774 4226
rect 471154 4102 471774 4170
rect 471154 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 471774 4102
rect 471154 3978 471774 4046
rect 471154 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 471774 3978
rect 471154 -160 471774 3922
rect 471154 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 471774 -160
rect 471154 -284 471774 -216
rect 471154 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 471774 -284
rect 471154 -408 471774 -340
rect 471154 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 471774 -408
rect 471154 -532 471774 -464
rect 471154 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 471774 -532
rect 471154 -1644 471774 -588
rect 474874 10350 475494 18186
rect 474874 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 475494 10350
rect 474874 10226 475494 10294
rect 474874 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 475494 10226
rect 474874 10102 475494 10170
rect 474874 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 475494 10102
rect 474874 9978 475494 10046
rect 474874 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 475494 9978
rect 474874 -1120 475494 9922
rect 474874 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 475494 -1120
rect 474874 -1244 475494 -1176
rect 474874 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 475494 -1244
rect 474874 -1368 475494 -1300
rect 474874 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 475494 -1368
rect 474874 -1492 475494 -1424
rect 474874 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 475494 -1492
rect 474874 -1644 475494 -1548
rect 489154 4350 489774 18186
rect 489154 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 489774 4350
rect 489154 4226 489774 4294
rect 489154 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 489774 4226
rect 489154 4102 489774 4170
rect 489154 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 489774 4102
rect 489154 3978 489774 4046
rect 489154 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 489774 3978
rect 489154 -160 489774 3922
rect 489154 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 489774 -160
rect 489154 -284 489774 -216
rect 489154 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 489774 -284
rect 489154 -408 489774 -340
rect 489154 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 489774 -408
rect 489154 -532 489774 -464
rect 489154 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 489774 -532
rect 489154 -1644 489774 -588
rect 492874 10350 493494 18186
rect 492874 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 493494 10350
rect 492874 10226 493494 10294
rect 492874 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 493494 10226
rect 492874 10102 493494 10170
rect 492874 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 493494 10102
rect 492874 9978 493494 10046
rect 492874 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 493494 9978
rect 492874 -1120 493494 9922
rect 492874 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 493494 -1120
rect 492874 -1244 493494 -1176
rect 492874 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 493494 -1244
rect 492874 -1368 493494 -1300
rect 492874 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 493494 -1368
rect 492874 -1492 493494 -1424
rect 492874 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 493494 -1492
rect 492874 -1644 493494 -1548
rect 507154 4350 507774 18186
rect 507154 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 507774 4350
rect 507154 4226 507774 4294
rect 507154 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 507774 4226
rect 507154 4102 507774 4170
rect 507154 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 507774 4102
rect 507154 3978 507774 4046
rect 507154 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 507774 3978
rect 507154 -160 507774 3922
rect 507154 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 507774 -160
rect 507154 -284 507774 -216
rect 507154 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 507774 -284
rect 507154 -408 507774 -340
rect 507154 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 507774 -408
rect 507154 -532 507774 -464
rect 507154 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 507774 -532
rect 507154 -1644 507774 -588
rect 510874 10350 511494 18186
rect 510874 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 511494 10350
rect 510874 10226 511494 10294
rect 510874 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 511494 10226
rect 510874 10102 511494 10170
rect 510874 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 511494 10102
rect 510874 9978 511494 10046
rect 510874 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 511494 9978
rect 510874 -1120 511494 9922
rect 510874 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 511494 -1120
rect 510874 -1244 511494 -1176
rect 510874 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 511494 -1244
rect 510874 -1368 511494 -1300
rect 510874 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 511494 -1368
rect 510874 -1492 511494 -1424
rect 510874 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 511494 -1492
rect 510874 -1644 511494 -1548
rect 525154 4350 525774 21922
rect 525154 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 525774 4350
rect 525154 4226 525774 4294
rect 525154 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 525774 4226
rect 525154 4102 525774 4170
rect 525154 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 525774 4102
rect 525154 3978 525774 4046
rect 525154 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 525774 3978
rect 525154 -160 525774 3922
rect 525154 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 525774 -160
rect 525154 -284 525774 -216
rect 525154 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 525774 -284
rect 525154 -408 525774 -340
rect 525154 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 525774 -408
rect 525154 -532 525774 -464
rect 525154 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 525774 -532
rect 525154 -1644 525774 -588
rect 528874 598172 529494 598268
rect 528874 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 529494 598172
rect 528874 598048 529494 598116
rect 528874 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 529494 598048
rect 528874 597924 529494 597992
rect 528874 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 529494 597924
rect 528874 597800 529494 597868
rect 528874 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 529494 597800
rect 528874 586350 529494 597744
rect 528874 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 529494 586350
rect 528874 586226 529494 586294
rect 528874 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 529494 586226
rect 528874 586102 529494 586170
rect 528874 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 529494 586102
rect 528874 585978 529494 586046
rect 528874 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 529494 585978
rect 528874 568350 529494 585922
rect 528874 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 529494 568350
rect 528874 568226 529494 568294
rect 528874 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 529494 568226
rect 528874 568102 529494 568170
rect 528874 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 529494 568102
rect 528874 567978 529494 568046
rect 528874 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 529494 567978
rect 528874 550350 529494 567922
rect 528874 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 529494 550350
rect 528874 550226 529494 550294
rect 528874 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 529494 550226
rect 528874 550102 529494 550170
rect 528874 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 529494 550102
rect 528874 549978 529494 550046
rect 528874 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 529494 549978
rect 528874 532350 529494 549922
rect 528874 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 529494 532350
rect 528874 532226 529494 532294
rect 528874 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 529494 532226
rect 528874 532102 529494 532170
rect 528874 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 529494 532102
rect 528874 531978 529494 532046
rect 528874 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 529494 531978
rect 528874 514350 529494 531922
rect 528874 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 529494 514350
rect 528874 514226 529494 514294
rect 528874 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 529494 514226
rect 528874 514102 529494 514170
rect 528874 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 529494 514102
rect 528874 513978 529494 514046
rect 528874 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 529494 513978
rect 528874 496350 529494 513922
rect 528874 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 529494 496350
rect 528874 496226 529494 496294
rect 528874 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 529494 496226
rect 528874 496102 529494 496170
rect 528874 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 529494 496102
rect 528874 495978 529494 496046
rect 528874 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 529494 495978
rect 528874 478350 529494 495922
rect 528874 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 529494 478350
rect 528874 478226 529494 478294
rect 528874 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 529494 478226
rect 528874 478102 529494 478170
rect 528874 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 529494 478102
rect 528874 477978 529494 478046
rect 528874 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 529494 477978
rect 528874 460350 529494 477922
rect 528874 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 529494 460350
rect 528874 460226 529494 460294
rect 528874 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 529494 460226
rect 528874 460102 529494 460170
rect 528874 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 529494 460102
rect 528874 459978 529494 460046
rect 528874 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 529494 459978
rect 528874 442350 529494 459922
rect 528874 442294 528970 442350
rect 529026 442294 529094 442350
rect 529150 442294 529218 442350
rect 529274 442294 529342 442350
rect 529398 442294 529494 442350
rect 528874 442226 529494 442294
rect 528874 442170 528970 442226
rect 529026 442170 529094 442226
rect 529150 442170 529218 442226
rect 529274 442170 529342 442226
rect 529398 442170 529494 442226
rect 528874 442102 529494 442170
rect 528874 442046 528970 442102
rect 529026 442046 529094 442102
rect 529150 442046 529218 442102
rect 529274 442046 529342 442102
rect 529398 442046 529494 442102
rect 528874 441978 529494 442046
rect 528874 441922 528970 441978
rect 529026 441922 529094 441978
rect 529150 441922 529218 441978
rect 529274 441922 529342 441978
rect 529398 441922 529494 441978
rect 528874 424350 529494 441922
rect 528874 424294 528970 424350
rect 529026 424294 529094 424350
rect 529150 424294 529218 424350
rect 529274 424294 529342 424350
rect 529398 424294 529494 424350
rect 528874 424226 529494 424294
rect 528874 424170 528970 424226
rect 529026 424170 529094 424226
rect 529150 424170 529218 424226
rect 529274 424170 529342 424226
rect 529398 424170 529494 424226
rect 528874 424102 529494 424170
rect 528874 424046 528970 424102
rect 529026 424046 529094 424102
rect 529150 424046 529218 424102
rect 529274 424046 529342 424102
rect 529398 424046 529494 424102
rect 528874 423978 529494 424046
rect 528874 423922 528970 423978
rect 529026 423922 529094 423978
rect 529150 423922 529218 423978
rect 529274 423922 529342 423978
rect 529398 423922 529494 423978
rect 528874 406350 529494 423922
rect 528874 406294 528970 406350
rect 529026 406294 529094 406350
rect 529150 406294 529218 406350
rect 529274 406294 529342 406350
rect 529398 406294 529494 406350
rect 528874 406226 529494 406294
rect 528874 406170 528970 406226
rect 529026 406170 529094 406226
rect 529150 406170 529218 406226
rect 529274 406170 529342 406226
rect 529398 406170 529494 406226
rect 528874 406102 529494 406170
rect 528874 406046 528970 406102
rect 529026 406046 529094 406102
rect 529150 406046 529218 406102
rect 529274 406046 529342 406102
rect 529398 406046 529494 406102
rect 528874 405978 529494 406046
rect 528874 405922 528970 405978
rect 529026 405922 529094 405978
rect 529150 405922 529218 405978
rect 529274 405922 529342 405978
rect 529398 405922 529494 405978
rect 528874 388350 529494 405922
rect 528874 388294 528970 388350
rect 529026 388294 529094 388350
rect 529150 388294 529218 388350
rect 529274 388294 529342 388350
rect 529398 388294 529494 388350
rect 528874 388226 529494 388294
rect 528874 388170 528970 388226
rect 529026 388170 529094 388226
rect 529150 388170 529218 388226
rect 529274 388170 529342 388226
rect 529398 388170 529494 388226
rect 528874 388102 529494 388170
rect 528874 388046 528970 388102
rect 529026 388046 529094 388102
rect 529150 388046 529218 388102
rect 529274 388046 529342 388102
rect 529398 388046 529494 388102
rect 528874 387978 529494 388046
rect 528874 387922 528970 387978
rect 529026 387922 529094 387978
rect 529150 387922 529218 387978
rect 529274 387922 529342 387978
rect 529398 387922 529494 387978
rect 528874 370350 529494 387922
rect 528874 370294 528970 370350
rect 529026 370294 529094 370350
rect 529150 370294 529218 370350
rect 529274 370294 529342 370350
rect 529398 370294 529494 370350
rect 528874 370226 529494 370294
rect 528874 370170 528970 370226
rect 529026 370170 529094 370226
rect 529150 370170 529218 370226
rect 529274 370170 529342 370226
rect 529398 370170 529494 370226
rect 528874 370102 529494 370170
rect 528874 370046 528970 370102
rect 529026 370046 529094 370102
rect 529150 370046 529218 370102
rect 529274 370046 529342 370102
rect 529398 370046 529494 370102
rect 528874 369978 529494 370046
rect 528874 369922 528970 369978
rect 529026 369922 529094 369978
rect 529150 369922 529218 369978
rect 529274 369922 529342 369978
rect 529398 369922 529494 369978
rect 528874 352350 529494 369922
rect 528874 352294 528970 352350
rect 529026 352294 529094 352350
rect 529150 352294 529218 352350
rect 529274 352294 529342 352350
rect 529398 352294 529494 352350
rect 528874 352226 529494 352294
rect 528874 352170 528970 352226
rect 529026 352170 529094 352226
rect 529150 352170 529218 352226
rect 529274 352170 529342 352226
rect 529398 352170 529494 352226
rect 528874 352102 529494 352170
rect 528874 352046 528970 352102
rect 529026 352046 529094 352102
rect 529150 352046 529218 352102
rect 529274 352046 529342 352102
rect 529398 352046 529494 352102
rect 528874 351978 529494 352046
rect 528874 351922 528970 351978
rect 529026 351922 529094 351978
rect 529150 351922 529218 351978
rect 529274 351922 529342 351978
rect 529398 351922 529494 351978
rect 528874 334350 529494 351922
rect 528874 334294 528970 334350
rect 529026 334294 529094 334350
rect 529150 334294 529218 334350
rect 529274 334294 529342 334350
rect 529398 334294 529494 334350
rect 528874 334226 529494 334294
rect 528874 334170 528970 334226
rect 529026 334170 529094 334226
rect 529150 334170 529218 334226
rect 529274 334170 529342 334226
rect 529398 334170 529494 334226
rect 528874 334102 529494 334170
rect 528874 334046 528970 334102
rect 529026 334046 529094 334102
rect 529150 334046 529218 334102
rect 529274 334046 529342 334102
rect 529398 334046 529494 334102
rect 528874 333978 529494 334046
rect 528874 333922 528970 333978
rect 529026 333922 529094 333978
rect 529150 333922 529218 333978
rect 529274 333922 529342 333978
rect 529398 333922 529494 333978
rect 528874 316350 529494 333922
rect 528874 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 529494 316350
rect 528874 316226 529494 316294
rect 528874 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 529494 316226
rect 528874 316102 529494 316170
rect 528874 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 529494 316102
rect 528874 315978 529494 316046
rect 528874 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 529494 315978
rect 528874 298350 529494 315922
rect 528874 298294 528970 298350
rect 529026 298294 529094 298350
rect 529150 298294 529218 298350
rect 529274 298294 529342 298350
rect 529398 298294 529494 298350
rect 528874 298226 529494 298294
rect 528874 298170 528970 298226
rect 529026 298170 529094 298226
rect 529150 298170 529218 298226
rect 529274 298170 529342 298226
rect 529398 298170 529494 298226
rect 528874 298102 529494 298170
rect 528874 298046 528970 298102
rect 529026 298046 529094 298102
rect 529150 298046 529218 298102
rect 529274 298046 529342 298102
rect 529398 298046 529494 298102
rect 528874 297978 529494 298046
rect 528874 297922 528970 297978
rect 529026 297922 529094 297978
rect 529150 297922 529218 297978
rect 529274 297922 529342 297978
rect 529398 297922 529494 297978
rect 528874 280350 529494 297922
rect 528874 280294 528970 280350
rect 529026 280294 529094 280350
rect 529150 280294 529218 280350
rect 529274 280294 529342 280350
rect 529398 280294 529494 280350
rect 528874 280226 529494 280294
rect 528874 280170 528970 280226
rect 529026 280170 529094 280226
rect 529150 280170 529218 280226
rect 529274 280170 529342 280226
rect 529398 280170 529494 280226
rect 528874 280102 529494 280170
rect 528874 280046 528970 280102
rect 529026 280046 529094 280102
rect 529150 280046 529218 280102
rect 529274 280046 529342 280102
rect 529398 280046 529494 280102
rect 528874 279978 529494 280046
rect 528874 279922 528970 279978
rect 529026 279922 529094 279978
rect 529150 279922 529218 279978
rect 529274 279922 529342 279978
rect 529398 279922 529494 279978
rect 528874 262350 529494 279922
rect 528874 262294 528970 262350
rect 529026 262294 529094 262350
rect 529150 262294 529218 262350
rect 529274 262294 529342 262350
rect 529398 262294 529494 262350
rect 528874 262226 529494 262294
rect 528874 262170 528970 262226
rect 529026 262170 529094 262226
rect 529150 262170 529218 262226
rect 529274 262170 529342 262226
rect 529398 262170 529494 262226
rect 528874 262102 529494 262170
rect 528874 262046 528970 262102
rect 529026 262046 529094 262102
rect 529150 262046 529218 262102
rect 529274 262046 529342 262102
rect 529398 262046 529494 262102
rect 528874 261978 529494 262046
rect 528874 261922 528970 261978
rect 529026 261922 529094 261978
rect 529150 261922 529218 261978
rect 529274 261922 529342 261978
rect 529398 261922 529494 261978
rect 528874 244350 529494 261922
rect 528874 244294 528970 244350
rect 529026 244294 529094 244350
rect 529150 244294 529218 244350
rect 529274 244294 529342 244350
rect 529398 244294 529494 244350
rect 528874 244226 529494 244294
rect 528874 244170 528970 244226
rect 529026 244170 529094 244226
rect 529150 244170 529218 244226
rect 529274 244170 529342 244226
rect 529398 244170 529494 244226
rect 528874 244102 529494 244170
rect 528874 244046 528970 244102
rect 529026 244046 529094 244102
rect 529150 244046 529218 244102
rect 529274 244046 529342 244102
rect 529398 244046 529494 244102
rect 528874 243978 529494 244046
rect 528874 243922 528970 243978
rect 529026 243922 529094 243978
rect 529150 243922 529218 243978
rect 529274 243922 529342 243978
rect 529398 243922 529494 243978
rect 528874 226350 529494 243922
rect 528874 226294 528970 226350
rect 529026 226294 529094 226350
rect 529150 226294 529218 226350
rect 529274 226294 529342 226350
rect 529398 226294 529494 226350
rect 528874 226226 529494 226294
rect 528874 226170 528970 226226
rect 529026 226170 529094 226226
rect 529150 226170 529218 226226
rect 529274 226170 529342 226226
rect 529398 226170 529494 226226
rect 528874 226102 529494 226170
rect 528874 226046 528970 226102
rect 529026 226046 529094 226102
rect 529150 226046 529218 226102
rect 529274 226046 529342 226102
rect 529398 226046 529494 226102
rect 528874 225978 529494 226046
rect 528874 225922 528970 225978
rect 529026 225922 529094 225978
rect 529150 225922 529218 225978
rect 529274 225922 529342 225978
rect 529398 225922 529494 225978
rect 528874 208350 529494 225922
rect 528874 208294 528970 208350
rect 529026 208294 529094 208350
rect 529150 208294 529218 208350
rect 529274 208294 529342 208350
rect 529398 208294 529494 208350
rect 528874 208226 529494 208294
rect 528874 208170 528970 208226
rect 529026 208170 529094 208226
rect 529150 208170 529218 208226
rect 529274 208170 529342 208226
rect 529398 208170 529494 208226
rect 528874 208102 529494 208170
rect 528874 208046 528970 208102
rect 529026 208046 529094 208102
rect 529150 208046 529218 208102
rect 529274 208046 529342 208102
rect 529398 208046 529494 208102
rect 528874 207978 529494 208046
rect 528874 207922 528970 207978
rect 529026 207922 529094 207978
rect 529150 207922 529218 207978
rect 529274 207922 529342 207978
rect 529398 207922 529494 207978
rect 528874 190350 529494 207922
rect 528874 190294 528970 190350
rect 529026 190294 529094 190350
rect 529150 190294 529218 190350
rect 529274 190294 529342 190350
rect 529398 190294 529494 190350
rect 528874 190226 529494 190294
rect 528874 190170 528970 190226
rect 529026 190170 529094 190226
rect 529150 190170 529218 190226
rect 529274 190170 529342 190226
rect 529398 190170 529494 190226
rect 528874 190102 529494 190170
rect 528874 190046 528970 190102
rect 529026 190046 529094 190102
rect 529150 190046 529218 190102
rect 529274 190046 529342 190102
rect 529398 190046 529494 190102
rect 528874 189978 529494 190046
rect 528874 189922 528970 189978
rect 529026 189922 529094 189978
rect 529150 189922 529218 189978
rect 529274 189922 529342 189978
rect 529398 189922 529494 189978
rect 528874 172350 529494 189922
rect 528874 172294 528970 172350
rect 529026 172294 529094 172350
rect 529150 172294 529218 172350
rect 529274 172294 529342 172350
rect 529398 172294 529494 172350
rect 528874 172226 529494 172294
rect 528874 172170 528970 172226
rect 529026 172170 529094 172226
rect 529150 172170 529218 172226
rect 529274 172170 529342 172226
rect 529398 172170 529494 172226
rect 528874 172102 529494 172170
rect 528874 172046 528970 172102
rect 529026 172046 529094 172102
rect 529150 172046 529218 172102
rect 529274 172046 529342 172102
rect 529398 172046 529494 172102
rect 528874 171978 529494 172046
rect 528874 171922 528970 171978
rect 529026 171922 529094 171978
rect 529150 171922 529218 171978
rect 529274 171922 529342 171978
rect 529398 171922 529494 171978
rect 528874 154350 529494 171922
rect 528874 154294 528970 154350
rect 529026 154294 529094 154350
rect 529150 154294 529218 154350
rect 529274 154294 529342 154350
rect 529398 154294 529494 154350
rect 528874 154226 529494 154294
rect 528874 154170 528970 154226
rect 529026 154170 529094 154226
rect 529150 154170 529218 154226
rect 529274 154170 529342 154226
rect 529398 154170 529494 154226
rect 528874 154102 529494 154170
rect 528874 154046 528970 154102
rect 529026 154046 529094 154102
rect 529150 154046 529218 154102
rect 529274 154046 529342 154102
rect 529398 154046 529494 154102
rect 528874 153978 529494 154046
rect 528874 153922 528970 153978
rect 529026 153922 529094 153978
rect 529150 153922 529218 153978
rect 529274 153922 529342 153978
rect 529398 153922 529494 153978
rect 528874 136350 529494 153922
rect 528874 136294 528970 136350
rect 529026 136294 529094 136350
rect 529150 136294 529218 136350
rect 529274 136294 529342 136350
rect 529398 136294 529494 136350
rect 528874 136226 529494 136294
rect 528874 136170 528970 136226
rect 529026 136170 529094 136226
rect 529150 136170 529218 136226
rect 529274 136170 529342 136226
rect 529398 136170 529494 136226
rect 528874 136102 529494 136170
rect 528874 136046 528970 136102
rect 529026 136046 529094 136102
rect 529150 136046 529218 136102
rect 529274 136046 529342 136102
rect 529398 136046 529494 136102
rect 528874 135978 529494 136046
rect 528874 135922 528970 135978
rect 529026 135922 529094 135978
rect 529150 135922 529218 135978
rect 529274 135922 529342 135978
rect 529398 135922 529494 135978
rect 528874 118350 529494 135922
rect 528874 118294 528970 118350
rect 529026 118294 529094 118350
rect 529150 118294 529218 118350
rect 529274 118294 529342 118350
rect 529398 118294 529494 118350
rect 528874 118226 529494 118294
rect 528874 118170 528970 118226
rect 529026 118170 529094 118226
rect 529150 118170 529218 118226
rect 529274 118170 529342 118226
rect 529398 118170 529494 118226
rect 528874 118102 529494 118170
rect 528874 118046 528970 118102
rect 529026 118046 529094 118102
rect 529150 118046 529218 118102
rect 529274 118046 529342 118102
rect 529398 118046 529494 118102
rect 528874 117978 529494 118046
rect 528874 117922 528970 117978
rect 529026 117922 529094 117978
rect 529150 117922 529218 117978
rect 529274 117922 529342 117978
rect 529398 117922 529494 117978
rect 528874 100350 529494 117922
rect 528874 100294 528970 100350
rect 529026 100294 529094 100350
rect 529150 100294 529218 100350
rect 529274 100294 529342 100350
rect 529398 100294 529494 100350
rect 528874 100226 529494 100294
rect 528874 100170 528970 100226
rect 529026 100170 529094 100226
rect 529150 100170 529218 100226
rect 529274 100170 529342 100226
rect 529398 100170 529494 100226
rect 528874 100102 529494 100170
rect 528874 100046 528970 100102
rect 529026 100046 529094 100102
rect 529150 100046 529218 100102
rect 529274 100046 529342 100102
rect 529398 100046 529494 100102
rect 528874 99978 529494 100046
rect 528874 99922 528970 99978
rect 529026 99922 529094 99978
rect 529150 99922 529218 99978
rect 529274 99922 529342 99978
rect 529398 99922 529494 99978
rect 528874 82350 529494 99922
rect 528874 82294 528970 82350
rect 529026 82294 529094 82350
rect 529150 82294 529218 82350
rect 529274 82294 529342 82350
rect 529398 82294 529494 82350
rect 528874 82226 529494 82294
rect 528874 82170 528970 82226
rect 529026 82170 529094 82226
rect 529150 82170 529218 82226
rect 529274 82170 529342 82226
rect 529398 82170 529494 82226
rect 528874 82102 529494 82170
rect 528874 82046 528970 82102
rect 529026 82046 529094 82102
rect 529150 82046 529218 82102
rect 529274 82046 529342 82102
rect 529398 82046 529494 82102
rect 528874 81978 529494 82046
rect 528874 81922 528970 81978
rect 529026 81922 529094 81978
rect 529150 81922 529218 81978
rect 529274 81922 529342 81978
rect 529398 81922 529494 81978
rect 528874 64350 529494 81922
rect 528874 64294 528970 64350
rect 529026 64294 529094 64350
rect 529150 64294 529218 64350
rect 529274 64294 529342 64350
rect 529398 64294 529494 64350
rect 528874 64226 529494 64294
rect 528874 64170 528970 64226
rect 529026 64170 529094 64226
rect 529150 64170 529218 64226
rect 529274 64170 529342 64226
rect 529398 64170 529494 64226
rect 528874 64102 529494 64170
rect 528874 64046 528970 64102
rect 529026 64046 529094 64102
rect 529150 64046 529218 64102
rect 529274 64046 529342 64102
rect 529398 64046 529494 64102
rect 528874 63978 529494 64046
rect 528874 63922 528970 63978
rect 529026 63922 529094 63978
rect 529150 63922 529218 63978
rect 529274 63922 529342 63978
rect 529398 63922 529494 63978
rect 528874 46350 529494 63922
rect 528874 46294 528970 46350
rect 529026 46294 529094 46350
rect 529150 46294 529218 46350
rect 529274 46294 529342 46350
rect 529398 46294 529494 46350
rect 528874 46226 529494 46294
rect 528874 46170 528970 46226
rect 529026 46170 529094 46226
rect 529150 46170 529218 46226
rect 529274 46170 529342 46226
rect 529398 46170 529494 46226
rect 528874 46102 529494 46170
rect 528874 46046 528970 46102
rect 529026 46046 529094 46102
rect 529150 46046 529218 46102
rect 529274 46046 529342 46102
rect 529398 46046 529494 46102
rect 528874 45978 529494 46046
rect 528874 45922 528970 45978
rect 529026 45922 529094 45978
rect 529150 45922 529218 45978
rect 529274 45922 529342 45978
rect 529398 45922 529494 45978
rect 528874 28350 529494 45922
rect 528874 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 529494 28350
rect 528874 28226 529494 28294
rect 528874 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 529494 28226
rect 528874 28102 529494 28170
rect 528874 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 529494 28102
rect 528874 27978 529494 28046
rect 528874 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 529494 27978
rect 528874 10350 529494 27922
rect 528874 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 529494 10350
rect 528874 10226 529494 10294
rect 528874 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 529494 10226
rect 528874 10102 529494 10170
rect 528874 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 529494 10102
rect 528874 9978 529494 10046
rect 528874 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 529494 9978
rect 528874 -1120 529494 9922
rect 528874 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 529494 -1120
rect 528874 -1244 529494 -1176
rect 528874 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 529494 -1244
rect 528874 -1368 529494 -1300
rect 528874 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 529494 -1368
rect 528874 -1492 529494 -1424
rect 528874 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 529494 -1492
rect 528874 -1644 529494 -1548
rect 543154 597212 543774 598268
rect 543154 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 543774 597212
rect 543154 597088 543774 597156
rect 543154 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 543774 597088
rect 543154 596964 543774 597032
rect 543154 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 543774 596964
rect 543154 596840 543774 596908
rect 543154 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 543774 596840
rect 543154 580350 543774 596784
rect 543154 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 543774 580350
rect 543154 580226 543774 580294
rect 543154 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 543774 580226
rect 543154 580102 543774 580170
rect 543154 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 543774 580102
rect 543154 579978 543774 580046
rect 543154 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 543774 579978
rect 543154 562350 543774 579922
rect 543154 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 543774 562350
rect 543154 562226 543774 562294
rect 543154 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 543774 562226
rect 543154 562102 543774 562170
rect 543154 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 543774 562102
rect 543154 561978 543774 562046
rect 543154 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 543774 561978
rect 543154 544350 543774 561922
rect 543154 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 543774 544350
rect 543154 544226 543774 544294
rect 543154 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 543774 544226
rect 543154 544102 543774 544170
rect 543154 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 543774 544102
rect 543154 543978 543774 544046
rect 543154 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 543774 543978
rect 543154 526350 543774 543922
rect 543154 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 543774 526350
rect 543154 526226 543774 526294
rect 543154 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 543774 526226
rect 543154 526102 543774 526170
rect 543154 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 543774 526102
rect 543154 525978 543774 526046
rect 543154 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 543774 525978
rect 543154 508350 543774 525922
rect 543154 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 543774 508350
rect 543154 508226 543774 508294
rect 543154 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 543774 508226
rect 543154 508102 543774 508170
rect 543154 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 543774 508102
rect 543154 507978 543774 508046
rect 543154 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 543774 507978
rect 543154 490350 543774 507922
rect 543154 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 543774 490350
rect 543154 490226 543774 490294
rect 543154 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 543774 490226
rect 543154 490102 543774 490170
rect 543154 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 543774 490102
rect 543154 489978 543774 490046
rect 543154 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 543774 489978
rect 543154 472350 543774 489922
rect 543154 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 543774 472350
rect 543154 472226 543774 472294
rect 543154 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 543774 472226
rect 543154 472102 543774 472170
rect 543154 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 543774 472102
rect 543154 471978 543774 472046
rect 543154 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 543774 471978
rect 543154 454350 543774 471922
rect 543154 454294 543250 454350
rect 543306 454294 543374 454350
rect 543430 454294 543498 454350
rect 543554 454294 543622 454350
rect 543678 454294 543774 454350
rect 543154 454226 543774 454294
rect 543154 454170 543250 454226
rect 543306 454170 543374 454226
rect 543430 454170 543498 454226
rect 543554 454170 543622 454226
rect 543678 454170 543774 454226
rect 543154 454102 543774 454170
rect 543154 454046 543250 454102
rect 543306 454046 543374 454102
rect 543430 454046 543498 454102
rect 543554 454046 543622 454102
rect 543678 454046 543774 454102
rect 543154 453978 543774 454046
rect 543154 453922 543250 453978
rect 543306 453922 543374 453978
rect 543430 453922 543498 453978
rect 543554 453922 543622 453978
rect 543678 453922 543774 453978
rect 543154 436350 543774 453922
rect 543154 436294 543250 436350
rect 543306 436294 543374 436350
rect 543430 436294 543498 436350
rect 543554 436294 543622 436350
rect 543678 436294 543774 436350
rect 543154 436226 543774 436294
rect 543154 436170 543250 436226
rect 543306 436170 543374 436226
rect 543430 436170 543498 436226
rect 543554 436170 543622 436226
rect 543678 436170 543774 436226
rect 543154 436102 543774 436170
rect 543154 436046 543250 436102
rect 543306 436046 543374 436102
rect 543430 436046 543498 436102
rect 543554 436046 543622 436102
rect 543678 436046 543774 436102
rect 543154 435978 543774 436046
rect 543154 435922 543250 435978
rect 543306 435922 543374 435978
rect 543430 435922 543498 435978
rect 543554 435922 543622 435978
rect 543678 435922 543774 435978
rect 543154 418350 543774 435922
rect 543154 418294 543250 418350
rect 543306 418294 543374 418350
rect 543430 418294 543498 418350
rect 543554 418294 543622 418350
rect 543678 418294 543774 418350
rect 543154 418226 543774 418294
rect 543154 418170 543250 418226
rect 543306 418170 543374 418226
rect 543430 418170 543498 418226
rect 543554 418170 543622 418226
rect 543678 418170 543774 418226
rect 543154 418102 543774 418170
rect 543154 418046 543250 418102
rect 543306 418046 543374 418102
rect 543430 418046 543498 418102
rect 543554 418046 543622 418102
rect 543678 418046 543774 418102
rect 543154 417978 543774 418046
rect 543154 417922 543250 417978
rect 543306 417922 543374 417978
rect 543430 417922 543498 417978
rect 543554 417922 543622 417978
rect 543678 417922 543774 417978
rect 543154 400350 543774 417922
rect 543154 400294 543250 400350
rect 543306 400294 543374 400350
rect 543430 400294 543498 400350
rect 543554 400294 543622 400350
rect 543678 400294 543774 400350
rect 543154 400226 543774 400294
rect 543154 400170 543250 400226
rect 543306 400170 543374 400226
rect 543430 400170 543498 400226
rect 543554 400170 543622 400226
rect 543678 400170 543774 400226
rect 543154 400102 543774 400170
rect 543154 400046 543250 400102
rect 543306 400046 543374 400102
rect 543430 400046 543498 400102
rect 543554 400046 543622 400102
rect 543678 400046 543774 400102
rect 543154 399978 543774 400046
rect 543154 399922 543250 399978
rect 543306 399922 543374 399978
rect 543430 399922 543498 399978
rect 543554 399922 543622 399978
rect 543678 399922 543774 399978
rect 543154 382350 543774 399922
rect 543154 382294 543250 382350
rect 543306 382294 543374 382350
rect 543430 382294 543498 382350
rect 543554 382294 543622 382350
rect 543678 382294 543774 382350
rect 543154 382226 543774 382294
rect 543154 382170 543250 382226
rect 543306 382170 543374 382226
rect 543430 382170 543498 382226
rect 543554 382170 543622 382226
rect 543678 382170 543774 382226
rect 543154 382102 543774 382170
rect 543154 382046 543250 382102
rect 543306 382046 543374 382102
rect 543430 382046 543498 382102
rect 543554 382046 543622 382102
rect 543678 382046 543774 382102
rect 543154 381978 543774 382046
rect 543154 381922 543250 381978
rect 543306 381922 543374 381978
rect 543430 381922 543498 381978
rect 543554 381922 543622 381978
rect 543678 381922 543774 381978
rect 543154 364350 543774 381922
rect 543154 364294 543250 364350
rect 543306 364294 543374 364350
rect 543430 364294 543498 364350
rect 543554 364294 543622 364350
rect 543678 364294 543774 364350
rect 543154 364226 543774 364294
rect 543154 364170 543250 364226
rect 543306 364170 543374 364226
rect 543430 364170 543498 364226
rect 543554 364170 543622 364226
rect 543678 364170 543774 364226
rect 543154 364102 543774 364170
rect 543154 364046 543250 364102
rect 543306 364046 543374 364102
rect 543430 364046 543498 364102
rect 543554 364046 543622 364102
rect 543678 364046 543774 364102
rect 543154 363978 543774 364046
rect 543154 363922 543250 363978
rect 543306 363922 543374 363978
rect 543430 363922 543498 363978
rect 543554 363922 543622 363978
rect 543678 363922 543774 363978
rect 543154 346350 543774 363922
rect 543154 346294 543250 346350
rect 543306 346294 543374 346350
rect 543430 346294 543498 346350
rect 543554 346294 543622 346350
rect 543678 346294 543774 346350
rect 543154 346226 543774 346294
rect 543154 346170 543250 346226
rect 543306 346170 543374 346226
rect 543430 346170 543498 346226
rect 543554 346170 543622 346226
rect 543678 346170 543774 346226
rect 543154 346102 543774 346170
rect 543154 346046 543250 346102
rect 543306 346046 543374 346102
rect 543430 346046 543498 346102
rect 543554 346046 543622 346102
rect 543678 346046 543774 346102
rect 543154 345978 543774 346046
rect 543154 345922 543250 345978
rect 543306 345922 543374 345978
rect 543430 345922 543498 345978
rect 543554 345922 543622 345978
rect 543678 345922 543774 345978
rect 543154 328350 543774 345922
rect 543154 328294 543250 328350
rect 543306 328294 543374 328350
rect 543430 328294 543498 328350
rect 543554 328294 543622 328350
rect 543678 328294 543774 328350
rect 543154 328226 543774 328294
rect 543154 328170 543250 328226
rect 543306 328170 543374 328226
rect 543430 328170 543498 328226
rect 543554 328170 543622 328226
rect 543678 328170 543774 328226
rect 543154 328102 543774 328170
rect 543154 328046 543250 328102
rect 543306 328046 543374 328102
rect 543430 328046 543498 328102
rect 543554 328046 543622 328102
rect 543678 328046 543774 328102
rect 543154 327978 543774 328046
rect 543154 327922 543250 327978
rect 543306 327922 543374 327978
rect 543430 327922 543498 327978
rect 543554 327922 543622 327978
rect 543678 327922 543774 327978
rect 543154 310350 543774 327922
rect 543154 310294 543250 310350
rect 543306 310294 543374 310350
rect 543430 310294 543498 310350
rect 543554 310294 543622 310350
rect 543678 310294 543774 310350
rect 543154 310226 543774 310294
rect 543154 310170 543250 310226
rect 543306 310170 543374 310226
rect 543430 310170 543498 310226
rect 543554 310170 543622 310226
rect 543678 310170 543774 310226
rect 543154 310102 543774 310170
rect 543154 310046 543250 310102
rect 543306 310046 543374 310102
rect 543430 310046 543498 310102
rect 543554 310046 543622 310102
rect 543678 310046 543774 310102
rect 543154 309978 543774 310046
rect 543154 309922 543250 309978
rect 543306 309922 543374 309978
rect 543430 309922 543498 309978
rect 543554 309922 543622 309978
rect 543678 309922 543774 309978
rect 543154 292350 543774 309922
rect 543154 292294 543250 292350
rect 543306 292294 543374 292350
rect 543430 292294 543498 292350
rect 543554 292294 543622 292350
rect 543678 292294 543774 292350
rect 543154 292226 543774 292294
rect 543154 292170 543250 292226
rect 543306 292170 543374 292226
rect 543430 292170 543498 292226
rect 543554 292170 543622 292226
rect 543678 292170 543774 292226
rect 543154 292102 543774 292170
rect 543154 292046 543250 292102
rect 543306 292046 543374 292102
rect 543430 292046 543498 292102
rect 543554 292046 543622 292102
rect 543678 292046 543774 292102
rect 543154 291978 543774 292046
rect 543154 291922 543250 291978
rect 543306 291922 543374 291978
rect 543430 291922 543498 291978
rect 543554 291922 543622 291978
rect 543678 291922 543774 291978
rect 543154 274350 543774 291922
rect 543154 274294 543250 274350
rect 543306 274294 543374 274350
rect 543430 274294 543498 274350
rect 543554 274294 543622 274350
rect 543678 274294 543774 274350
rect 543154 274226 543774 274294
rect 543154 274170 543250 274226
rect 543306 274170 543374 274226
rect 543430 274170 543498 274226
rect 543554 274170 543622 274226
rect 543678 274170 543774 274226
rect 543154 274102 543774 274170
rect 543154 274046 543250 274102
rect 543306 274046 543374 274102
rect 543430 274046 543498 274102
rect 543554 274046 543622 274102
rect 543678 274046 543774 274102
rect 543154 273978 543774 274046
rect 543154 273922 543250 273978
rect 543306 273922 543374 273978
rect 543430 273922 543498 273978
rect 543554 273922 543622 273978
rect 543678 273922 543774 273978
rect 543154 256350 543774 273922
rect 543154 256294 543250 256350
rect 543306 256294 543374 256350
rect 543430 256294 543498 256350
rect 543554 256294 543622 256350
rect 543678 256294 543774 256350
rect 543154 256226 543774 256294
rect 543154 256170 543250 256226
rect 543306 256170 543374 256226
rect 543430 256170 543498 256226
rect 543554 256170 543622 256226
rect 543678 256170 543774 256226
rect 543154 256102 543774 256170
rect 543154 256046 543250 256102
rect 543306 256046 543374 256102
rect 543430 256046 543498 256102
rect 543554 256046 543622 256102
rect 543678 256046 543774 256102
rect 543154 255978 543774 256046
rect 543154 255922 543250 255978
rect 543306 255922 543374 255978
rect 543430 255922 543498 255978
rect 543554 255922 543622 255978
rect 543678 255922 543774 255978
rect 543154 238350 543774 255922
rect 543154 238294 543250 238350
rect 543306 238294 543374 238350
rect 543430 238294 543498 238350
rect 543554 238294 543622 238350
rect 543678 238294 543774 238350
rect 543154 238226 543774 238294
rect 543154 238170 543250 238226
rect 543306 238170 543374 238226
rect 543430 238170 543498 238226
rect 543554 238170 543622 238226
rect 543678 238170 543774 238226
rect 543154 238102 543774 238170
rect 543154 238046 543250 238102
rect 543306 238046 543374 238102
rect 543430 238046 543498 238102
rect 543554 238046 543622 238102
rect 543678 238046 543774 238102
rect 543154 237978 543774 238046
rect 543154 237922 543250 237978
rect 543306 237922 543374 237978
rect 543430 237922 543498 237978
rect 543554 237922 543622 237978
rect 543678 237922 543774 237978
rect 543154 220350 543774 237922
rect 543154 220294 543250 220350
rect 543306 220294 543374 220350
rect 543430 220294 543498 220350
rect 543554 220294 543622 220350
rect 543678 220294 543774 220350
rect 543154 220226 543774 220294
rect 543154 220170 543250 220226
rect 543306 220170 543374 220226
rect 543430 220170 543498 220226
rect 543554 220170 543622 220226
rect 543678 220170 543774 220226
rect 543154 220102 543774 220170
rect 543154 220046 543250 220102
rect 543306 220046 543374 220102
rect 543430 220046 543498 220102
rect 543554 220046 543622 220102
rect 543678 220046 543774 220102
rect 543154 219978 543774 220046
rect 543154 219922 543250 219978
rect 543306 219922 543374 219978
rect 543430 219922 543498 219978
rect 543554 219922 543622 219978
rect 543678 219922 543774 219978
rect 543154 202350 543774 219922
rect 543154 202294 543250 202350
rect 543306 202294 543374 202350
rect 543430 202294 543498 202350
rect 543554 202294 543622 202350
rect 543678 202294 543774 202350
rect 543154 202226 543774 202294
rect 543154 202170 543250 202226
rect 543306 202170 543374 202226
rect 543430 202170 543498 202226
rect 543554 202170 543622 202226
rect 543678 202170 543774 202226
rect 543154 202102 543774 202170
rect 543154 202046 543250 202102
rect 543306 202046 543374 202102
rect 543430 202046 543498 202102
rect 543554 202046 543622 202102
rect 543678 202046 543774 202102
rect 543154 201978 543774 202046
rect 543154 201922 543250 201978
rect 543306 201922 543374 201978
rect 543430 201922 543498 201978
rect 543554 201922 543622 201978
rect 543678 201922 543774 201978
rect 543154 184350 543774 201922
rect 543154 184294 543250 184350
rect 543306 184294 543374 184350
rect 543430 184294 543498 184350
rect 543554 184294 543622 184350
rect 543678 184294 543774 184350
rect 543154 184226 543774 184294
rect 543154 184170 543250 184226
rect 543306 184170 543374 184226
rect 543430 184170 543498 184226
rect 543554 184170 543622 184226
rect 543678 184170 543774 184226
rect 543154 184102 543774 184170
rect 543154 184046 543250 184102
rect 543306 184046 543374 184102
rect 543430 184046 543498 184102
rect 543554 184046 543622 184102
rect 543678 184046 543774 184102
rect 543154 183978 543774 184046
rect 543154 183922 543250 183978
rect 543306 183922 543374 183978
rect 543430 183922 543498 183978
rect 543554 183922 543622 183978
rect 543678 183922 543774 183978
rect 543154 166350 543774 183922
rect 543154 166294 543250 166350
rect 543306 166294 543374 166350
rect 543430 166294 543498 166350
rect 543554 166294 543622 166350
rect 543678 166294 543774 166350
rect 543154 166226 543774 166294
rect 543154 166170 543250 166226
rect 543306 166170 543374 166226
rect 543430 166170 543498 166226
rect 543554 166170 543622 166226
rect 543678 166170 543774 166226
rect 543154 166102 543774 166170
rect 543154 166046 543250 166102
rect 543306 166046 543374 166102
rect 543430 166046 543498 166102
rect 543554 166046 543622 166102
rect 543678 166046 543774 166102
rect 543154 165978 543774 166046
rect 543154 165922 543250 165978
rect 543306 165922 543374 165978
rect 543430 165922 543498 165978
rect 543554 165922 543622 165978
rect 543678 165922 543774 165978
rect 543154 148350 543774 165922
rect 543154 148294 543250 148350
rect 543306 148294 543374 148350
rect 543430 148294 543498 148350
rect 543554 148294 543622 148350
rect 543678 148294 543774 148350
rect 543154 148226 543774 148294
rect 543154 148170 543250 148226
rect 543306 148170 543374 148226
rect 543430 148170 543498 148226
rect 543554 148170 543622 148226
rect 543678 148170 543774 148226
rect 543154 148102 543774 148170
rect 543154 148046 543250 148102
rect 543306 148046 543374 148102
rect 543430 148046 543498 148102
rect 543554 148046 543622 148102
rect 543678 148046 543774 148102
rect 543154 147978 543774 148046
rect 543154 147922 543250 147978
rect 543306 147922 543374 147978
rect 543430 147922 543498 147978
rect 543554 147922 543622 147978
rect 543678 147922 543774 147978
rect 543154 130350 543774 147922
rect 543154 130294 543250 130350
rect 543306 130294 543374 130350
rect 543430 130294 543498 130350
rect 543554 130294 543622 130350
rect 543678 130294 543774 130350
rect 543154 130226 543774 130294
rect 543154 130170 543250 130226
rect 543306 130170 543374 130226
rect 543430 130170 543498 130226
rect 543554 130170 543622 130226
rect 543678 130170 543774 130226
rect 543154 130102 543774 130170
rect 543154 130046 543250 130102
rect 543306 130046 543374 130102
rect 543430 130046 543498 130102
rect 543554 130046 543622 130102
rect 543678 130046 543774 130102
rect 543154 129978 543774 130046
rect 543154 129922 543250 129978
rect 543306 129922 543374 129978
rect 543430 129922 543498 129978
rect 543554 129922 543622 129978
rect 543678 129922 543774 129978
rect 543154 112350 543774 129922
rect 543154 112294 543250 112350
rect 543306 112294 543374 112350
rect 543430 112294 543498 112350
rect 543554 112294 543622 112350
rect 543678 112294 543774 112350
rect 543154 112226 543774 112294
rect 543154 112170 543250 112226
rect 543306 112170 543374 112226
rect 543430 112170 543498 112226
rect 543554 112170 543622 112226
rect 543678 112170 543774 112226
rect 543154 112102 543774 112170
rect 543154 112046 543250 112102
rect 543306 112046 543374 112102
rect 543430 112046 543498 112102
rect 543554 112046 543622 112102
rect 543678 112046 543774 112102
rect 543154 111978 543774 112046
rect 543154 111922 543250 111978
rect 543306 111922 543374 111978
rect 543430 111922 543498 111978
rect 543554 111922 543622 111978
rect 543678 111922 543774 111978
rect 543154 94350 543774 111922
rect 543154 94294 543250 94350
rect 543306 94294 543374 94350
rect 543430 94294 543498 94350
rect 543554 94294 543622 94350
rect 543678 94294 543774 94350
rect 543154 94226 543774 94294
rect 543154 94170 543250 94226
rect 543306 94170 543374 94226
rect 543430 94170 543498 94226
rect 543554 94170 543622 94226
rect 543678 94170 543774 94226
rect 543154 94102 543774 94170
rect 543154 94046 543250 94102
rect 543306 94046 543374 94102
rect 543430 94046 543498 94102
rect 543554 94046 543622 94102
rect 543678 94046 543774 94102
rect 543154 93978 543774 94046
rect 543154 93922 543250 93978
rect 543306 93922 543374 93978
rect 543430 93922 543498 93978
rect 543554 93922 543622 93978
rect 543678 93922 543774 93978
rect 543154 76350 543774 93922
rect 543154 76294 543250 76350
rect 543306 76294 543374 76350
rect 543430 76294 543498 76350
rect 543554 76294 543622 76350
rect 543678 76294 543774 76350
rect 543154 76226 543774 76294
rect 543154 76170 543250 76226
rect 543306 76170 543374 76226
rect 543430 76170 543498 76226
rect 543554 76170 543622 76226
rect 543678 76170 543774 76226
rect 543154 76102 543774 76170
rect 543154 76046 543250 76102
rect 543306 76046 543374 76102
rect 543430 76046 543498 76102
rect 543554 76046 543622 76102
rect 543678 76046 543774 76102
rect 543154 75978 543774 76046
rect 543154 75922 543250 75978
rect 543306 75922 543374 75978
rect 543430 75922 543498 75978
rect 543554 75922 543622 75978
rect 543678 75922 543774 75978
rect 543154 58350 543774 75922
rect 543154 58294 543250 58350
rect 543306 58294 543374 58350
rect 543430 58294 543498 58350
rect 543554 58294 543622 58350
rect 543678 58294 543774 58350
rect 543154 58226 543774 58294
rect 543154 58170 543250 58226
rect 543306 58170 543374 58226
rect 543430 58170 543498 58226
rect 543554 58170 543622 58226
rect 543678 58170 543774 58226
rect 543154 58102 543774 58170
rect 543154 58046 543250 58102
rect 543306 58046 543374 58102
rect 543430 58046 543498 58102
rect 543554 58046 543622 58102
rect 543678 58046 543774 58102
rect 543154 57978 543774 58046
rect 543154 57922 543250 57978
rect 543306 57922 543374 57978
rect 543430 57922 543498 57978
rect 543554 57922 543622 57978
rect 543678 57922 543774 57978
rect 543154 40350 543774 57922
rect 543154 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 543774 40350
rect 543154 40226 543774 40294
rect 543154 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 543774 40226
rect 543154 40102 543774 40170
rect 543154 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 543774 40102
rect 543154 39978 543774 40046
rect 543154 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 543774 39978
rect 543154 22350 543774 39922
rect 543154 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 543774 22350
rect 543154 22226 543774 22294
rect 543154 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 543774 22226
rect 543154 22102 543774 22170
rect 543154 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 543774 22102
rect 543154 21978 543774 22046
rect 543154 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 543774 21978
rect 543154 4350 543774 21922
rect 543154 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 543774 4350
rect 543154 4226 543774 4294
rect 543154 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 543774 4226
rect 543154 4102 543774 4170
rect 543154 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 543774 4102
rect 543154 3978 543774 4046
rect 543154 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 543774 3978
rect 543154 -160 543774 3922
rect 543154 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 543774 -160
rect 543154 -284 543774 -216
rect 543154 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 543774 -284
rect 543154 -408 543774 -340
rect 543154 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 543774 -408
rect 543154 -532 543774 -464
rect 543154 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 543774 -532
rect 543154 -1644 543774 -588
rect 546874 598172 547494 598268
rect 546874 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 547494 598172
rect 546874 598048 547494 598116
rect 546874 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 547494 598048
rect 546874 597924 547494 597992
rect 546874 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 547494 597924
rect 546874 597800 547494 597868
rect 546874 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 547494 597800
rect 546874 586350 547494 597744
rect 546874 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 547494 586350
rect 546874 586226 547494 586294
rect 546874 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 547494 586226
rect 546874 586102 547494 586170
rect 546874 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 547494 586102
rect 546874 585978 547494 586046
rect 546874 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 547494 585978
rect 546874 568350 547494 585922
rect 546874 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 547494 568350
rect 546874 568226 547494 568294
rect 546874 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 547494 568226
rect 546874 568102 547494 568170
rect 546874 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 547494 568102
rect 546874 567978 547494 568046
rect 546874 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 547494 567978
rect 546874 550350 547494 567922
rect 546874 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 547494 550350
rect 546874 550226 547494 550294
rect 546874 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 547494 550226
rect 546874 550102 547494 550170
rect 546874 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 547494 550102
rect 546874 549978 547494 550046
rect 546874 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 547494 549978
rect 546874 532350 547494 549922
rect 546874 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 547494 532350
rect 546874 532226 547494 532294
rect 546874 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 547494 532226
rect 546874 532102 547494 532170
rect 546874 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 547494 532102
rect 546874 531978 547494 532046
rect 546874 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 547494 531978
rect 546874 514350 547494 531922
rect 546874 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 547494 514350
rect 546874 514226 547494 514294
rect 546874 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 547494 514226
rect 546874 514102 547494 514170
rect 546874 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 547494 514102
rect 546874 513978 547494 514046
rect 546874 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 547494 513978
rect 546874 496350 547494 513922
rect 546874 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 547494 496350
rect 546874 496226 547494 496294
rect 546874 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 547494 496226
rect 546874 496102 547494 496170
rect 546874 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 547494 496102
rect 546874 495978 547494 496046
rect 546874 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 547494 495978
rect 546874 478350 547494 495922
rect 546874 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 547494 478350
rect 546874 478226 547494 478294
rect 546874 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 547494 478226
rect 546874 478102 547494 478170
rect 546874 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 547494 478102
rect 546874 477978 547494 478046
rect 546874 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 547494 477978
rect 546874 460350 547494 477922
rect 546874 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 547494 460350
rect 546874 460226 547494 460294
rect 546874 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 547494 460226
rect 546874 460102 547494 460170
rect 546874 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 547494 460102
rect 546874 459978 547494 460046
rect 546874 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 547494 459978
rect 546874 442350 547494 459922
rect 546874 442294 546970 442350
rect 547026 442294 547094 442350
rect 547150 442294 547218 442350
rect 547274 442294 547342 442350
rect 547398 442294 547494 442350
rect 546874 442226 547494 442294
rect 546874 442170 546970 442226
rect 547026 442170 547094 442226
rect 547150 442170 547218 442226
rect 547274 442170 547342 442226
rect 547398 442170 547494 442226
rect 546874 442102 547494 442170
rect 546874 442046 546970 442102
rect 547026 442046 547094 442102
rect 547150 442046 547218 442102
rect 547274 442046 547342 442102
rect 547398 442046 547494 442102
rect 546874 441978 547494 442046
rect 546874 441922 546970 441978
rect 547026 441922 547094 441978
rect 547150 441922 547218 441978
rect 547274 441922 547342 441978
rect 547398 441922 547494 441978
rect 546874 424350 547494 441922
rect 546874 424294 546970 424350
rect 547026 424294 547094 424350
rect 547150 424294 547218 424350
rect 547274 424294 547342 424350
rect 547398 424294 547494 424350
rect 546874 424226 547494 424294
rect 546874 424170 546970 424226
rect 547026 424170 547094 424226
rect 547150 424170 547218 424226
rect 547274 424170 547342 424226
rect 547398 424170 547494 424226
rect 546874 424102 547494 424170
rect 546874 424046 546970 424102
rect 547026 424046 547094 424102
rect 547150 424046 547218 424102
rect 547274 424046 547342 424102
rect 547398 424046 547494 424102
rect 546874 423978 547494 424046
rect 546874 423922 546970 423978
rect 547026 423922 547094 423978
rect 547150 423922 547218 423978
rect 547274 423922 547342 423978
rect 547398 423922 547494 423978
rect 546874 406350 547494 423922
rect 546874 406294 546970 406350
rect 547026 406294 547094 406350
rect 547150 406294 547218 406350
rect 547274 406294 547342 406350
rect 547398 406294 547494 406350
rect 546874 406226 547494 406294
rect 546874 406170 546970 406226
rect 547026 406170 547094 406226
rect 547150 406170 547218 406226
rect 547274 406170 547342 406226
rect 547398 406170 547494 406226
rect 546874 406102 547494 406170
rect 546874 406046 546970 406102
rect 547026 406046 547094 406102
rect 547150 406046 547218 406102
rect 547274 406046 547342 406102
rect 547398 406046 547494 406102
rect 546874 405978 547494 406046
rect 546874 405922 546970 405978
rect 547026 405922 547094 405978
rect 547150 405922 547218 405978
rect 547274 405922 547342 405978
rect 547398 405922 547494 405978
rect 546874 388350 547494 405922
rect 546874 388294 546970 388350
rect 547026 388294 547094 388350
rect 547150 388294 547218 388350
rect 547274 388294 547342 388350
rect 547398 388294 547494 388350
rect 546874 388226 547494 388294
rect 546874 388170 546970 388226
rect 547026 388170 547094 388226
rect 547150 388170 547218 388226
rect 547274 388170 547342 388226
rect 547398 388170 547494 388226
rect 546874 388102 547494 388170
rect 546874 388046 546970 388102
rect 547026 388046 547094 388102
rect 547150 388046 547218 388102
rect 547274 388046 547342 388102
rect 547398 388046 547494 388102
rect 546874 387978 547494 388046
rect 546874 387922 546970 387978
rect 547026 387922 547094 387978
rect 547150 387922 547218 387978
rect 547274 387922 547342 387978
rect 547398 387922 547494 387978
rect 546874 370350 547494 387922
rect 546874 370294 546970 370350
rect 547026 370294 547094 370350
rect 547150 370294 547218 370350
rect 547274 370294 547342 370350
rect 547398 370294 547494 370350
rect 546874 370226 547494 370294
rect 546874 370170 546970 370226
rect 547026 370170 547094 370226
rect 547150 370170 547218 370226
rect 547274 370170 547342 370226
rect 547398 370170 547494 370226
rect 546874 370102 547494 370170
rect 546874 370046 546970 370102
rect 547026 370046 547094 370102
rect 547150 370046 547218 370102
rect 547274 370046 547342 370102
rect 547398 370046 547494 370102
rect 546874 369978 547494 370046
rect 546874 369922 546970 369978
rect 547026 369922 547094 369978
rect 547150 369922 547218 369978
rect 547274 369922 547342 369978
rect 547398 369922 547494 369978
rect 546874 352350 547494 369922
rect 546874 352294 546970 352350
rect 547026 352294 547094 352350
rect 547150 352294 547218 352350
rect 547274 352294 547342 352350
rect 547398 352294 547494 352350
rect 546874 352226 547494 352294
rect 546874 352170 546970 352226
rect 547026 352170 547094 352226
rect 547150 352170 547218 352226
rect 547274 352170 547342 352226
rect 547398 352170 547494 352226
rect 546874 352102 547494 352170
rect 546874 352046 546970 352102
rect 547026 352046 547094 352102
rect 547150 352046 547218 352102
rect 547274 352046 547342 352102
rect 547398 352046 547494 352102
rect 546874 351978 547494 352046
rect 546874 351922 546970 351978
rect 547026 351922 547094 351978
rect 547150 351922 547218 351978
rect 547274 351922 547342 351978
rect 547398 351922 547494 351978
rect 546874 334350 547494 351922
rect 546874 334294 546970 334350
rect 547026 334294 547094 334350
rect 547150 334294 547218 334350
rect 547274 334294 547342 334350
rect 547398 334294 547494 334350
rect 546874 334226 547494 334294
rect 546874 334170 546970 334226
rect 547026 334170 547094 334226
rect 547150 334170 547218 334226
rect 547274 334170 547342 334226
rect 547398 334170 547494 334226
rect 546874 334102 547494 334170
rect 546874 334046 546970 334102
rect 547026 334046 547094 334102
rect 547150 334046 547218 334102
rect 547274 334046 547342 334102
rect 547398 334046 547494 334102
rect 546874 333978 547494 334046
rect 546874 333922 546970 333978
rect 547026 333922 547094 333978
rect 547150 333922 547218 333978
rect 547274 333922 547342 333978
rect 547398 333922 547494 333978
rect 546874 316350 547494 333922
rect 546874 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 547494 316350
rect 546874 316226 547494 316294
rect 546874 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 547494 316226
rect 546874 316102 547494 316170
rect 546874 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 547494 316102
rect 546874 315978 547494 316046
rect 546874 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 547494 315978
rect 546874 298350 547494 315922
rect 546874 298294 546970 298350
rect 547026 298294 547094 298350
rect 547150 298294 547218 298350
rect 547274 298294 547342 298350
rect 547398 298294 547494 298350
rect 546874 298226 547494 298294
rect 546874 298170 546970 298226
rect 547026 298170 547094 298226
rect 547150 298170 547218 298226
rect 547274 298170 547342 298226
rect 547398 298170 547494 298226
rect 546874 298102 547494 298170
rect 546874 298046 546970 298102
rect 547026 298046 547094 298102
rect 547150 298046 547218 298102
rect 547274 298046 547342 298102
rect 547398 298046 547494 298102
rect 546874 297978 547494 298046
rect 546874 297922 546970 297978
rect 547026 297922 547094 297978
rect 547150 297922 547218 297978
rect 547274 297922 547342 297978
rect 547398 297922 547494 297978
rect 546874 280350 547494 297922
rect 546874 280294 546970 280350
rect 547026 280294 547094 280350
rect 547150 280294 547218 280350
rect 547274 280294 547342 280350
rect 547398 280294 547494 280350
rect 546874 280226 547494 280294
rect 546874 280170 546970 280226
rect 547026 280170 547094 280226
rect 547150 280170 547218 280226
rect 547274 280170 547342 280226
rect 547398 280170 547494 280226
rect 546874 280102 547494 280170
rect 546874 280046 546970 280102
rect 547026 280046 547094 280102
rect 547150 280046 547218 280102
rect 547274 280046 547342 280102
rect 547398 280046 547494 280102
rect 546874 279978 547494 280046
rect 546874 279922 546970 279978
rect 547026 279922 547094 279978
rect 547150 279922 547218 279978
rect 547274 279922 547342 279978
rect 547398 279922 547494 279978
rect 546874 262350 547494 279922
rect 546874 262294 546970 262350
rect 547026 262294 547094 262350
rect 547150 262294 547218 262350
rect 547274 262294 547342 262350
rect 547398 262294 547494 262350
rect 546874 262226 547494 262294
rect 546874 262170 546970 262226
rect 547026 262170 547094 262226
rect 547150 262170 547218 262226
rect 547274 262170 547342 262226
rect 547398 262170 547494 262226
rect 546874 262102 547494 262170
rect 546874 262046 546970 262102
rect 547026 262046 547094 262102
rect 547150 262046 547218 262102
rect 547274 262046 547342 262102
rect 547398 262046 547494 262102
rect 546874 261978 547494 262046
rect 546874 261922 546970 261978
rect 547026 261922 547094 261978
rect 547150 261922 547218 261978
rect 547274 261922 547342 261978
rect 547398 261922 547494 261978
rect 546874 244350 547494 261922
rect 546874 244294 546970 244350
rect 547026 244294 547094 244350
rect 547150 244294 547218 244350
rect 547274 244294 547342 244350
rect 547398 244294 547494 244350
rect 546874 244226 547494 244294
rect 546874 244170 546970 244226
rect 547026 244170 547094 244226
rect 547150 244170 547218 244226
rect 547274 244170 547342 244226
rect 547398 244170 547494 244226
rect 546874 244102 547494 244170
rect 546874 244046 546970 244102
rect 547026 244046 547094 244102
rect 547150 244046 547218 244102
rect 547274 244046 547342 244102
rect 547398 244046 547494 244102
rect 546874 243978 547494 244046
rect 546874 243922 546970 243978
rect 547026 243922 547094 243978
rect 547150 243922 547218 243978
rect 547274 243922 547342 243978
rect 547398 243922 547494 243978
rect 546874 226350 547494 243922
rect 546874 226294 546970 226350
rect 547026 226294 547094 226350
rect 547150 226294 547218 226350
rect 547274 226294 547342 226350
rect 547398 226294 547494 226350
rect 546874 226226 547494 226294
rect 546874 226170 546970 226226
rect 547026 226170 547094 226226
rect 547150 226170 547218 226226
rect 547274 226170 547342 226226
rect 547398 226170 547494 226226
rect 546874 226102 547494 226170
rect 546874 226046 546970 226102
rect 547026 226046 547094 226102
rect 547150 226046 547218 226102
rect 547274 226046 547342 226102
rect 547398 226046 547494 226102
rect 546874 225978 547494 226046
rect 546874 225922 546970 225978
rect 547026 225922 547094 225978
rect 547150 225922 547218 225978
rect 547274 225922 547342 225978
rect 547398 225922 547494 225978
rect 546874 208350 547494 225922
rect 546874 208294 546970 208350
rect 547026 208294 547094 208350
rect 547150 208294 547218 208350
rect 547274 208294 547342 208350
rect 547398 208294 547494 208350
rect 546874 208226 547494 208294
rect 546874 208170 546970 208226
rect 547026 208170 547094 208226
rect 547150 208170 547218 208226
rect 547274 208170 547342 208226
rect 547398 208170 547494 208226
rect 546874 208102 547494 208170
rect 546874 208046 546970 208102
rect 547026 208046 547094 208102
rect 547150 208046 547218 208102
rect 547274 208046 547342 208102
rect 547398 208046 547494 208102
rect 546874 207978 547494 208046
rect 546874 207922 546970 207978
rect 547026 207922 547094 207978
rect 547150 207922 547218 207978
rect 547274 207922 547342 207978
rect 547398 207922 547494 207978
rect 546874 190350 547494 207922
rect 546874 190294 546970 190350
rect 547026 190294 547094 190350
rect 547150 190294 547218 190350
rect 547274 190294 547342 190350
rect 547398 190294 547494 190350
rect 546874 190226 547494 190294
rect 546874 190170 546970 190226
rect 547026 190170 547094 190226
rect 547150 190170 547218 190226
rect 547274 190170 547342 190226
rect 547398 190170 547494 190226
rect 546874 190102 547494 190170
rect 546874 190046 546970 190102
rect 547026 190046 547094 190102
rect 547150 190046 547218 190102
rect 547274 190046 547342 190102
rect 547398 190046 547494 190102
rect 546874 189978 547494 190046
rect 546874 189922 546970 189978
rect 547026 189922 547094 189978
rect 547150 189922 547218 189978
rect 547274 189922 547342 189978
rect 547398 189922 547494 189978
rect 546874 172350 547494 189922
rect 546874 172294 546970 172350
rect 547026 172294 547094 172350
rect 547150 172294 547218 172350
rect 547274 172294 547342 172350
rect 547398 172294 547494 172350
rect 546874 172226 547494 172294
rect 546874 172170 546970 172226
rect 547026 172170 547094 172226
rect 547150 172170 547218 172226
rect 547274 172170 547342 172226
rect 547398 172170 547494 172226
rect 546874 172102 547494 172170
rect 546874 172046 546970 172102
rect 547026 172046 547094 172102
rect 547150 172046 547218 172102
rect 547274 172046 547342 172102
rect 547398 172046 547494 172102
rect 546874 171978 547494 172046
rect 546874 171922 546970 171978
rect 547026 171922 547094 171978
rect 547150 171922 547218 171978
rect 547274 171922 547342 171978
rect 547398 171922 547494 171978
rect 546874 154350 547494 171922
rect 546874 154294 546970 154350
rect 547026 154294 547094 154350
rect 547150 154294 547218 154350
rect 547274 154294 547342 154350
rect 547398 154294 547494 154350
rect 546874 154226 547494 154294
rect 546874 154170 546970 154226
rect 547026 154170 547094 154226
rect 547150 154170 547218 154226
rect 547274 154170 547342 154226
rect 547398 154170 547494 154226
rect 546874 154102 547494 154170
rect 546874 154046 546970 154102
rect 547026 154046 547094 154102
rect 547150 154046 547218 154102
rect 547274 154046 547342 154102
rect 547398 154046 547494 154102
rect 546874 153978 547494 154046
rect 546874 153922 546970 153978
rect 547026 153922 547094 153978
rect 547150 153922 547218 153978
rect 547274 153922 547342 153978
rect 547398 153922 547494 153978
rect 546874 136350 547494 153922
rect 546874 136294 546970 136350
rect 547026 136294 547094 136350
rect 547150 136294 547218 136350
rect 547274 136294 547342 136350
rect 547398 136294 547494 136350
rect 546874 136226 547494 136294
rect 546874 136170 546970 136226
rect 547026 136170 547094 136226
rect 547150 136170 547218 136226
rect 547274 136170 547342 136226
rect 547398 136170 547494 136226
rect 546874 136102 547494 136170
rect 546874 136046 546970 136102
rect 547026 136046 547094 136102
rect 547150 136046 547218 136102
rect 547274 136046 547342 136102
rect 547398 136046 547494 136102
rect 546874 135978 547494 136046
rect 546874 135922 546970 135978
rect 547026 135922 547094 135978
rect 547150 135922 547218 135978
rect 547274 135922 547342 135978
rect 547398 135922 547494 135978
rect 546874 118350 547494 135922
rect 546874 118294 546970 118350
rect 547026 118294 547094 118350
rect 547150 118294 547218 118350
rect 547274 118294 547342 118350
rect 547398 118294 547494 118350
rect 546874 118226 547494 118294
rect 546874 118170 546970 118226
rect 547026 118170 547094 118226
rect 547150 118170 547218 118226
rect 547274 118170 547342 118226
rect 547398 118170 547494 118226
rect 546874 118102 547494 118170
rect 546874 118046 546970 118102
rect 547026 118046 547094 118102
rect 547150 118046 547218 118102
rect 547274 118046 547342 118102
rect 547398 118046 547494 118102
rect 546874 117978 547494 118046
rect 546874 117922 546970 117978
rect 547026 117922 547094 117978
rect 547150 117922 547218 117978
rect 547274 117922 547342 117978
rect 547398 117922 547494 117978
rect 546874 100350 547494 117922
rect 546874 100294 546970 100350
rect 547026 100294 547094 100350
rect 547150 100294 547218 100350
rect 547274 100294 547342 100350
rect 547398 100294 547494 100350
rect 546874 100226 547494 100294
rect 546874 100170 546970 100226
rect 547026 100170 547094 100226
rect 547150 100170 547218 100226
rect 547274 100170 547342 100226
rect 547398 100170 547494 100226
rect 546874 100102 547494 100170
rect 546874 100046 546970 100102
rect 547026 100046 547094 100102
rect 547150 100046 547218 100102
rect 547274 100046 547342 100102
rect 547398 100046 547494 100102
rect 546874 99978 547494 100046
rect 546874 99922 546970 99978
rect 547026 99922 547094 99978
rect 547150 99922 547218 99978
rect 547274 99922 547342 99978
rect 547398 99922 547494 99978
rect 546874 82350 547494 99922
rect 546874 82294 546970 82350
rect 547026 82294 547094 82350
rect 547150 82294 547218 82350
rect 547274 82294 547342 82350
rect 547398 82294 547494 82350
rect 546874 82226 547494 82294
rect 546874 82170 546970 82226
rect 547026 82170 547094 82226
rect 547150 82170 547218 82226
rect 547274 82170 547342 82226
rect 547398 82170 547494 82226
rect 546874 82102 547494 82170
rect 546874 82046 546970 82102
rect 547026 82046 547094 82102
rect 547150 82046 547218 82102
rect 547274 82046 547342 82102
rect 547398 82046 547494 82102
rect 546874 81978 547494 82046
rect 546874 81922 546970 81978
rect 547026 81922 547094 81978
rect 547150 81922 547218 81978
rect 547274 81922 547342 81978
rect 547398 81922 547494 81978
rect 546874 64350 547494 81922
rect 546874 64294 546970 64350
rect 547026 64294 547094 64350
rect 547150 64294 547218 64350
rect 547274 64294 547342 64350
rect 547398 64294 547494 64350
rect 546874 64226 547494 64294
rect 546874 64170 546970 64226
rect 547026 64170 547094 64226
rect 547150 64170 547218 64226
rect 547274 64170 547342 64226
rect 547398 64170 547494 64226
rect 546874 64102 547494 64170
rect 546874 64046 546970 64102
rect 547026 64046 547094 64102
rect 547150 64046 547218 64102
rect 547274 64046 547342 64102
rect 547398 64046 547494 64102
rect 546874 63978 547494 64046
rect 546874 63922 546970 63978
rect 547026 63922 547094 63978
rect 547150 63922 547218 63978
rect 547274 63922 547342 63978
rect 547398 63922 547494 63978
rect 546874 46350 547494 63922
rect 546874 46294 546970 46350
rect 547026 46294 547094 46350
rect 547150 46294 547218 46350
rect 547274 46294 547342 46350
rect 547398 46294 547494 46350
rect 546874 46226 547494 46294
rect 546874 46170 546970 46226
rect 547026 46170 547094 46226
rect 547150 46170 547218 46226
rect 547274 46170 547342 46226
rect 547398 46170 547494 46226
rect 546874 46102 547494 46170
rect 546874 46046 546970 46102
rect 547026 46046 547094 46102
rect 547150 46046 547218 46102
rect 547274 46046 547342 46102
rect 547398 46046 547494 46102
rect 546874 45978 547494 46046
rect 546874 45922 546970 45978
rect 547026 45922 547094 45978
rect 547150 45922 547218 45978
rect 547274 45922 547342 45978
rect 547398 45922 547494 45978
rect 546874 28350 547494 45922
rect 546874 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 547494 28350
rect 546874 28226 547494 28294
rect 546874 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 547494 28226
rect 546874 28102 547494 28170
rect 546874 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 547494 28102
rect 546874 27978 547494 28046
rect 546874 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 547494 27978
rect 546874 10350 547494 27922
rect 546874 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 547494 10350
rect 546874 10226 547494 10294
rect 546874 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 547494 10226
rect 546874 10102 547494 10170
rect 546874 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 547494 10102
rect 546874 9978 547494 10046
rect 546874 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 547494 9978
rect 546874 -1120 547494 9922
rect 546874 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 547494 -1120
rect 546874 -1244 547494 -1176
rect 546874 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 547494 -1244
rect 546874 -1368 547494 -1300
rect 546874 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 547494 -1368
rect 546874 -1492 547494 -1424
rect 546874 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 547494 -1492
rect 546874 -1644 547494 -1548
rect 561154 597212 561774 598268
rect 561154 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 561774 597212
rect 561154 597088 561774 597156
rect 561154 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 561774 597088
rect 561154 596964 561774 597032
rect 561154 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 561774 596964
rect 561154 596840 561774 596908
rect 561154 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 561774 596840
rect 561154 580350 561774 596784
rect 561154 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 561774 580350
rect 561154 580226 561774 580294
rect 561154 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 561774 580226
rect 561154 580102 561774 580170
rect 561154 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 561774 580102
rect 561154 579978 561774 580046
rect 561154 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 561774 579978
rect 561154 562350 561774 579922
rect 561154 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 561774 562350
rect 561154 562226 561774 562294
rect 561154 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 561774 562226
rect 561154 562102 561774 562170
rect 561154 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 561774 562102
rect 561154 561978 561774 562046
rect 561154 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 561774 561978
rect 561154 544350 561774 561922
rect 561154 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 561774 544350
rect 561154 544226 561774 544294
rect 561154 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 561774 544226
rect 561154 544102 561774 544170
rect 561154 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 561774 544102
rect 561154 543978 561774 544046
rect 561154 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 561774 543978
rect 561154 526350 561774 543922
rect 561154 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 561774 526350
rect 561154 526226 561774 526294
rect 561154 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 561774 526226
rect 561154 526102 561774 526170
rect 561154 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 561774 526102
rect 561154 525978 561774 526046
rect 561154 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 561774 525978
rect 561154 508350 561774 525922
rect 561154 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 561774 508350
rect 561154 508226 561774 508294
rect 561154 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 561774 508226
rect 561154 508102 561774 508170
rect 561154 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 561774 508102
rect 561154 507978 561774 508046
rect 561154 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 561774 507978
rect 561154 490350 561774 507922
rect 561154 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 561774 490350
rect 561154 490226 561774 490294
rect 561154 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 561774 490226
rect 561154 490102 561774 490170
rect 561154 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 561774 490102
rect 561154 489978 561774 490046
rect 561154 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 561774 489978
rect 561154 472350 561774 489922
rect 561154 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 561774 472350
rect 561154 472226 561774 472294
rect 561154 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 561774 472226
rect 561154 472102 561774 472170
rect 561154 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 561774 472102
rect 561154 471978 561774 472046
rect 561154 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 561774 471978
rect 561154 454350 561774 471922
rect 561154 454294 561250 454350
rect 561306 454294 561374 454350
rect 561430 454294 561498 454350
rect 561554 454294 561622 454350
rect 561678 454294 561774 454350
rect 561154 454226 561774 454294
rect 561154 454170 561250 454226
rect 561306 454170 561374 454226
rect 561430 454170 561498 454226
rect 561554 454170 561622 454226
rect 561678 454170 561774 454226
rect 561154 454102 561774 454170
rect 561154 454046 561250 454102
rect 561306 454046 561374 454102
rect 561430 454046 561498 454102
rect 561554 454046 561622 454102
rect 561678 454046 561774 454102
rect 561154 453978 561774 454046
rect 561154 453922 561250 453978
rect 561306 453922 561374 453978
rect 561430 453922 561498 453978
rect 561554 453922 561622 453978
rect 561678 453922 561774 453978
rect 561154 436350 561774 453922
rect 561154 436294 561250 436350
rect 561306 436294 561374 436350
rect 561430 436294 561498 436350
rect 561554 436294 561622 436350
rect 561678 436294 561774 436350
rect 561154 436226 561774 436294
rect 561154 436170 561250 436226
rect 561306 436170 561374 436226
rect 561430 436170 561498 436226
rect 561554 436170 561622 436226
rect 561678 436170 561774 436226
rect 561154 436102 561774 436170
rect 561154 436046 561250 436102
rect 561306 436046 561374 436102
rect 561430 436046 561498 436102
rect 561554 436046 561622 436102
rect 561678 436046 561774 436102
rect 561154 435978 561774 436046
rect 561154 435922 561250 435978
rect 561306 435922 561374 435978
rect 561430 435922 561498 435978
rect 561554 435922 561622 435978
rect 561678 435922 561774 435978
rect 561154 418350 561774 435922
rect 561154 418294 561250 418350
rect 561306 418294 561374 418350
rect 561430 418294 561498 418350
rect 561554 418294 561622 418350
rect 561678 418294 561774 418350
rect 561154 418226 561774 418294
rect 561154 418170 561250 418226
rect 561306 418170 561374 418226
rect 561430 418170 561498 418226
rect 561554 418170 561622 418226
rect 561678 418170 561774 418226
rect 561154 418102 561774 418170
rect 561154 418046 561250 418102
rect 561306 418046 561374 418102
rect 561430 418046 561498 418102
rect 561554 418046 561622 418102
rect 561678 418046 561774 418102
rect 561154 417978 561774 418046
rect 561154 417922 561250 417978
rect 561306 417922 561374 417978
rect 561430 417922 561498 417978
rect 561554 417922 561622 417978
rect 561678 417922 561774 417978
rect 561154 400350 561774 417922
rect 561154 400294 561250 400350
rect 561306 400294 561374 400350
rect 561430 400294 561498 400350
rect 561554 400294 561622 400350
rect 561678 400294 561774 400350
rect 561154 400226 561774 400294
rect 561154 400170 561250 400226
rect 561306 400170 561374 400226
rect 561430 400170 561498 400226
rect 561554 400170 561622 400226
rect 561678 400170 561774 400226
rect 561154 400102 561774 400170
rect 561154 400046 561250 400102
rect 561306 400046 561374 400102
rect 561430 400046 561498 400102
rect 561554 400046 561622 400102
rect 561678 400046 561774 400102
rect 561154 399978 561774 400046
rect 561154 399922 561250 399978
rect 561306 399922 561374 399978
rect 561430 399922 561498 399978
rect 561554 399922 561622 399978
rect 561678 399922 561774 399978
rect 561154 382350 561774 399922
rect 561154 382294 561250 382350
rect 561306 382294 561374 382350
rect 561430 382294 561498 382350
rect 561554 382294 561622 382350
rect 561678 382294 561774 382350
rect 561154 382226 561774 382294
rect 561154 382170 561250 382226
rect 561306 382170 561374 382226
rect 561430 382170 561498 382226
rect 561554 382170 561622 382226
rect 561678 382170 561774 382226
rect 561154 382102 561774 382170
rect 561154 382046 561250 382102
rect 561306 382046 561374 382102
rect 561430 382046 561498 382102
rect 561554 382046 561622 382102
rect 561678 382046 561774 382102
rect 561154 381978 561774 382046
rect 561154 381922 561250 381978
rect 561306 381922 561374 381978
rect 561430 381922 561498 381978
rect 561554 381922 561622 381978
rect 561678 381922 561774 381978
rect 561154 364350 561774 381922
rect 561154 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 561774 364350
rect 561154 364226 561774 364294
rect 561154 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 561774 364226
rect 561154 364102 561774 364170
rect 561154 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 561774 364102
rect 561154 363978 561774 364046
rect 561154 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 561774 363978
rect 561154 346350 561774 363922
rect 561154 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 561774 346350
rect 561154 346226 561774 346294
rect 561154 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 561774 346226
rect 561154 346102 561774 346170
rect 561154 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 561774 346102
rect 561154 345978 561774 346046
rect 561154 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 561774 345978
rect 561154 328350 561774 345922
rect 561154 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 561774 328350
rect 561154 328226 561774 328294
rect 561154 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 561774 328226
rect 561154 328102 561774 328170
rect 561154 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 561774 328102
rect 561154 327978 561774 328046
rect 561154 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 561774 327978
rect 561154 310350 561774 327922
rect 561154 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 561774 310350
rect 561154 310226 561774 310294
rect 561154 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 561774 310226
rect 561154 310102 561774 310170
rect 561154 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 561774 310102
rect 561154 309978 561774 310046
rect 561154 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 561774 309978
rect 561154 292350 561774 309922
rect 561154 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 561774 292350
rect 561154 292226 561774 292294
rect 561154 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 561774 292226
rect 561154 292102 561774 292170
rect 561154 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 561774 292102
rect 561154 291978 561774 292046
rect 561154 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 561774 291978
rect 561154 274350 561774 291922
rect 561154 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 561774 274350
rect 561154 274226 561774 274294
rect 561154 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 561774 274226
rect 561154 274102 561774 274170
rect 561154 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 561774 274102
rect 561154 273978 561774 274046
rect 561154 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 561774 273978
rect 561154 256350 561774 273922
rect 561154 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 561774 256350
rect 561154 256226 561774 256294
rect 561154 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 561774 256226
rect 561154 256102 561774 256170
rect 561154 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 561774 256102
rect 561154 255978 561774 256046
rect 561154 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 561774 255978
rect 561154 238350 561774 255922
rect 561154 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 561774 238350
rect 561154 238226 561774 238294
rect 561154 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 561774 238226
rect 561154 238102 561774 238170
rect 561154 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 561774 238102
rect 561154 237978 561774 238046
rect 561154 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 561774 237978
rect 561154 220350 561774 237922
rect 561154 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 561774 220350
rect 561154 220226 561774 220294
rect 561154 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 561774 220226
rect 561154 220102 561774 220170
rect 561154 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 561774 220102
rect 561154 219978 561774 220046
rect 561154 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 561774 219978
rect 561154 202350 561774 219922
rect 561154 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 561774 202350
rect 561154 202226 561774 202294
rect 561154 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 561774 202226
rect 561154 202102 561774 202170
rect 561154 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 561774 202102
rect 561154 201978 561774 202046
rect 561154 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 561774 201978
rect 561154 184350 561774 201922
rect 561154 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 561774 184350
rect 561154 184226 561774 184294
rect 561154 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 561774 184226
rect 561154 184102 561774 184170
rect 561154 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 561774 184102
rect 561154 183978 561774 184046
rect 561154 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 561774 183978
rect 561154 166350 561774 183922
rect 561154 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 561774 166350
rect 561154 166226 561774 166294
rect 561154 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 561774 166226
rect 561154 166102 561774 166170
rect 561154 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 561774 166102
rect 561154 165978 561774 166046
rect 561154 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 561774 165978
rect 561154 148350 561774 165922
rect 561154 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 561774 148350
rect 561154 148226 561774 148294
rect 561154 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 561774 148226
rect 561154 148102 561774 148170
rect 561154 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 561774 148102
rect 561154 147978 561774 148046
rect 561154 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 561774 147978
rect 561154 130350 561774 147922
rect 561154 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 561774 130350
rect 561154 130226 561774 130294
rect 561154 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 561774 130226
rect 561154 130102 561774 130170
rect 561154 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 561774 130102
rect 561154 129978 561774 130046
rect 561154 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 561774 129978
rect 561154 112350 561774 129922
rect 561154 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 561774 112350
rect 561154 112226 561774 112294
rect 561154 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 561774 112226
rect 561154 112102 561774 112170
rect 561154 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 561774 112102
rect 561154 111978 561774 112046
rect 561154 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 561774 111978
rect 561154 94350 561774 111922
rect 561154 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 561774 94350
rect 561154 94226 561774 94294
rect 561154 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 561774 94226
rect 561154 94102 561774 94170
rect 561154 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 561774 94102
rect 561154 93978 561774 94046
rect 561154 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 561774 93978
rect 561154 76350 561774 93922
rect 561154 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 561774 76350
rect 561154 76226 561774 76294
rect 561154 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 561774 76226
rect 561154 76102 561774 76170
rect 561154 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 561774 76102
rect 561154 75978 561774 76046
rect 561154 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 561774 75978
rect 561154 58350 561774 75922
rect 561154 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 561774 58350
rect 561154 58226 561774 58294
rect 561154 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 561774 58226
rect 561154 58102 561774 58170
rect 561154 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 561774 58102
rect 561154 57978 561774 58046
rect 561154 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 561774 57978
rect 561154 40350 561774 57922
rect 561154 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 561774 40350
rect 561154 40226 561774 40294
rect 561154 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 561774 40226
rect 561154 40102 561774 40170
rect 561154 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 561774 40102
rect 561154 39978 561774 40046
rect 561154 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 561774 39978
rect 561154 22350 561774 39922
rect 561154 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 561774 22350
rect 561154 22226 561774 22294
rect 561154 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 561774 22226
rect 561154 22102 561774 22170
rect 561154 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 561774 22102
rect 561154 21978 561774 22046
rect 561154 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 561774 21978
rect 561154 4350 561774 21922
rect 561154 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 561774 4350
rect 561154 4226 561774 4294
rect 561154 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 561774 4226
rect 561154 4102 561774 4170
rect 561154 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 561774 4102
rect 561154 3978 561774 4046
rect 561154 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 561774 3978
rect 561154 -160 561774 3922
rect 561154 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 561774 -160
rect 561154 -284 561774 -216
rect 561154 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 561774 -284
rect 561154 -408 561774 -340
rect 561154 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 561774 -408
rect 561154 -532 561774 -464
rect 561154 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 561774 -532
rect 561154 -1644 561774 -588
rect 564874 598172 565494 598268
rect 564874 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 565494 598172
rect 564874 598048 565494 598116
rect 564874 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 565494 598048
rect 564874 597924 565494 597992
rect 564874 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 565494 597924
rect 564874 597800 565494 597868
rect 564874 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 565494 597800
rect 564874 586350 565494 597744
rect 564874 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 565494 586350
rect 564874 586226 565494 586294
rect 564874 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 565494 586226
rect 564874 586102 565494 586170
rect 564874 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 565494 586102
rect 564874 585978 565494 586046
rect 564874 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 565494 585978
rect 564874 568350 565494 585922
rect 564874 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 565494 568350
rect 564874 568226 565494 568294
rect 564874 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 565494 568226
rect 564874 568102 565494 568170
rect 564874 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 565494 568102
rect 564874 567978 565494 568046
rect 564874 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 565494 567978
rect 564874 550350 565494 567922
rect 564874 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 565494 550350
rect 564874 550226 565494 550294
rect 564874 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 565494 550226
rect 564874 550102 565494 550170
rect 564874 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 565494 550102
rect 564874 549978 565494 550046
rect 564874 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 565494 549978
rect 564874 532350 565494 549922
rect 564874 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 565494 532350
rect 564874 532226 565494 532294
rect 564874 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 565494 532226
rect 564874 532102 565494 532170
rect 564874 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 565494 532102
rect 564874 531978 565494 532046
rect 564874 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 565494 531978
rect 564874 514350 565494 531922
rect 564874 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 565494 514350
rect 564874 514226 565494 514294
rect 564874 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 565494 514226
rect 564874 514102 565494 514170
rect 564874 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 565494 514102
rect 564874 513978 565494 514046
rect 564874 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 565494 513978
rect 564874 496350 565494 513922
rect 564874 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 565494 496350
rect 564874 496226 565494 496294
rect 564874 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 565494 496226
rect 564874 496102 565494 496170
rect 564874 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 565494 496102
rect 564874 495978 565494 496046
rect 564874 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 565494 495978
rect 564874 478350 565494 495922
rect 564874 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 565494 478350
rect 564874 478226 565494 478294
rect 564874 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 565494 478226
rect 564874 478102 565494 478170
rect 564874 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 565494 478102
rect 564874 477978 565494 478046
rect 564874 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 565494 477978
rect 564874 460350 565494 477922
rect 564874 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 565494 460350
rect 564874 460226 565494 460294
rect 564874 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 565494 460226
rect 564874 460102 565494 460170
rect 564874 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 565494 460102
rect 564874 459978 565494 460046
rect 564874 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 565494 459978
rect 564874 442350 565494 459922
rect 564874 442294 564970 442350
rect 565026 442294 565094 442350
rect 565150 442294 565218 442350
rect 565274 442294 565342 442350
rect 565398 442294 565494 442350
rect 564874 442226 565494 442294
rect 564874 442170 564970 442226
rect 565026 442170 565094 442226
rect 565150 442170 565218 442226
rect 565274 442170 565342 442226
rect 565398 442170 565494 442226
rect 564874 442102 565494 442170
rect 564874 442046 564970 442102
rect 565026 442046 565094 442102
rect 565150 442046 565218 442102
rect 565274 442046 565342 442102
rect 565398 442046 565494 442102
rect 564874 441978 565494 442046
rect 564874 441922 564970 441978
rect 565026 441922 565094 441978
rect 565150 441922 565218 441978
rect 565274 441922 565342 441978
rect 565398 441922 565494 441978
rect 564874 424350 565494 441922
rect 564874 424294 564970 424350
rect 565026 424294 565094 424350
rect 565150 424294 565218 424350
rect 565274 424294 565342 424350
rect 565398 424294 565494 424350
rect 564874 424226 565494 424294
rect 564874 424170 564970 424226
rect 565026 424170 565094 424226
rect 565150 424170 565218 424226
rect 565274 424170 565342 424226
rect 565398 424170 565494 424226
rect 564874 424102 565494 424170
rect 564874 424046 564970 424102
rect 565026 424046 565094 424102
rect 565150 424046 565218 424102
rect 565274 424046 565342 424102
rect 565398 424046 565494 424102
rect 564874 423978 565494 424046
rect 564874 423922 564970 423978
rect 565026 423922 565094 423978
rect 565150 423922 565218 423978
rect 565274 423922 565342 423978
rect 565398 423922 565494 423978
rect 564874 406350 565494 423922
rect 564874 406294 564970 406350
rect 565026 406294 565094 406350
rect 565150 406294 565218 406350
rect 565274 406294 565342 406350
rect 565398 406294 565494 406350
rect 564874 406226 565494 406294
rect 564874 406170 564970 406226
rect 565026 406170 565094 406226
rect 565150 406170 565218 406226
rect 565274 406170 565342 406226
rect 565398 406170 565494 406226
rect 564874 406102 565494 406170
rect 564874 406046 564970 406102
rect 565026 406046 565094 406102
rect 565150 406046 565218 406102
rect 565274 406046 565342 406102
rect 565398 406046 565494 406102
rect 564874 405978 565494 406046
rect 564874 405922 564970 405978
rect 565026 405922 565094 405978
rect 565150 405922 565218 405978
rect 565274 405922 565342 405978
rect 565398 405922 565494 405978
rect 564874 388350 565494 405922
rect 564874 388294 564970 388350
rect 565026 388294 565094 388350
rect 565150 388294 565218 388350
rect 565274 388294 565342 388350
rect 565398 388294 565494 388350
rect 564874 388226 565494 388294
rect 564874 388170 564970 388226
rect 565026 388170 565094 388226
rect 565150 388170 565218 388226
rect 565274 388170 565342 388226
rect 565398 388170 565494 388226
rect 564874 388102 565494 388170
rect 564874 388046 564970 388102
rect 565026 388046 565094 388102
rect 565150 388046 565218 388102
rect 565274 388046 565342 388102
rect 565398 388046 565494 388102
rect 564874 387978 565494 388046
rect 564874 387922 564970 387978
rect 565026 387922 565094 387978
rect 565150 387922 565218 387978
rect 565274 387922 565342 387978
rect 565398 387922 565494 387978
rect 564874 370350 565494 387922
rect 564874 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 565494 370350
rect 564874 370226 565494 370294
rect 564874 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 565494 370226
rect 564874 370102 565494 370170
rect 564874 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 565494 370102
rect 564874 369978 565494 370046
rect 564874 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 565494 369978
rect 564874 352350 565494 369922
rect 564874 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 565494 352350
rect 564874 352226 565494 352294
rect 564874 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 565494 352226
rect 564874 352102 565494 352170
rect 564874 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 565494 352102
rect 564874 351978 565494 352046
rect 564874 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 565494 351978
rect 564874 334350 565494 351922
rect 564874 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 565494 334350
rect 564874 334226 565494 334294
rect 564874 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 565494 334226
rect 564874 334102 565494 334170
rect 564874 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 565494 334102
rect 564874 333978 565494 334046
rect 564874 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 565494 333978
rect 564874 316350 565494 333922
rect 564874 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 565494 316350
rect 564874 316226 565494 316294
rect 564874 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 565494 316226
rect 564874 316102 565494 316170
rect 564874 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 565494 316102
rect 564874 315978 565494 316046
rect 564874 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 565494 315978
rect 564874 298350 565494 315922
rect 564874 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 565494 298350
rect 564874 298226 565494 298294
rect 564874 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 565494 298226
rect 564874 298102 565494 298170
rect 564874 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 565494 298102
rect 564874 297978 565494 298046
rect 564874 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 565494 297978
rect 564874 280350 565494 297922
rect 564874 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 565494 280350
rect 564874 280226 565494 280294
rect 564874 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 565494 280226
rect 564874 280102 565494 280170
rect 564874 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 565494 280102
rect 564874 279978 565494 280046
rect 564874 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 565494 279978
rect 564874 262350 565494 279922
rect 564874 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 565494 262350
rect 564874 262226 565494 262294
rect 564874 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 565494 262226
rect 564874 262102 565494 262170
rect 564874 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 565494 262102
rect 564874 261978 565494 262046
rect 564874 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 565494 261978
rect 564874 244350 565494 261922
rect 564874 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 565494 244350
rect 564874 244226 565494 244294
rect 564874 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 565494 244226
rect 564874 244102 565494 244170
rect 564874 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 565494 244102
rect 564874 243978 565494 244046
rect 564874 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 565494 243978
rect 564874 226350 565494 243922
rect 564874 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 565494 226350
rect 564874 226226 565494 226294
rect 564874 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 565494 226226
rect 564874 226102 565494 226170
rect 564874 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 565494 226102
rect 564874 225978 565494 226046
rect 564874 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 565494 225978
rect 564874 208350 565494 225922
rect 564874 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 565494 208350
rect 564874 208226 565494 208294
rect 564874 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 565494 208226
rect 564874 208102 565494 208170
rect 564874 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 565494 208102
rect 564874 207978 565494 208046
rect 564874 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 565494 207978
rect 564874 190350 565494 207922
rect 564874 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 565494 190350
rect 564874 190226 565494 190294
rect 564874 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 565494 190226
rect 564874 190102 565494 190170
rect 564874 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 565494 190102
rect 564874 189978 565494 190046
rect 564874 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 565494 189978
rect 564874 172350 565494 189922
rect 564874 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 565494 172350
rect 564874 172226 565494 172294
rect 564874 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 565494 172226
rect 564874 172102 565494 172170
rect 564874 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 565494 172102
rect 564874 171978 565494 172046
rect 564874 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 565494 171978
rect 564874 154350 565494 171922
rect 564874 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 565494 154350
rect 564874 154226 565494 154294
rect 564874 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 565494 154226
rect 564874 154102 565494 154170
rect 564874 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 565494 154102
rect 564874 153978 565494 154046
rect 564874 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 565494 153978
rect 564874 136350 565494 153922
rect 564874 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 565494 136350
rect 564874 136226 565494 136294
rect 564874 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 565494 136226
rect 564874 136102 565494 136170
rect 564874 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 565494 136102
rect 564874 135978 565494 136046
rect 564874 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 565494 135978
rect 564874 118350 565494 135922
rect 564874 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 565494 118350
rect 564874 118226 565494 118294
rect 564874 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 565494 118226
rect 564874 118102 565494 118170
rect 564874 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 565494 118102
rect 564874 117978 565494 118046
rect 564874 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 565494 117978
rect 564874 100350 565494 117922
rect 564874 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 565494 100350
rect 564874 100226 565494 100294
rect 564874 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 565494 100226
rect 564874 100102 565494 100170
rect 564874 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 565494 100102
rect 564874 99978 565494 100046
rect 564874 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 565494 99978
rect 564874 82350 565494 99922
rect 564874 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 565494 82350
rect 564874 82226 565494 82294
rect 564874 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 565494 82226
rect 564874 82102 565494 82170
rect 564874 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 565494 82102
rect 564874 81978 565494 82046
rect 564874 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 565494 81978
rect 564874 64350 565494 81922
rect 564874 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 565494 64350
rect 564874 64226 565494 64294
rect 564874 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 565494 64226
rect 564874 64102 565494 64170
rect 564874 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 565494 64102
rect 564874 63978 565494 64046
rect 564874 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 565494 63978
rect 564874 46350 565494 63922
rect 564874 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 565494 46350
rect 564874 46226 565494 46294
rect 564874 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 565494 46226
rect 564874 46102 565494 46170
rect 564874 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 565494 46102
rect 564874 45978 565494 46046
rect 564874 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 565494 45978
rect 564874 28350 565494 45922
rect 564874 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 565494 28350
rect 564874 28226 565494 28294
rect 564874 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 565494 28226
rect 564874 28102 565494 28170
rect 564874 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 565494 28102
rect 564874 27978 565494 28046
rect 564874 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 565494 27978
rect 564874 10350 565494 27922
rect 564874 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 565494 10350
rect 564874 10226 565494 10294
rect 564874 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 565494 10226
rect 564874 10102 565494 10170
rect 564874 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 565494 10102
rect 564874 9978 565494 10046
rect 564874 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 565494 9978
rect 564874 -1120 565494 9922
rect 564874 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 565494 -1120
rect 564874 -1244 565494 -1176
rect 564874 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 565494 -1244
rect 564874 -1368 565494 -1300
rect 564874 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 565494 -1368
rect 564874 -1492 565494 -1424
rect 564874 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 565494 -1492
rect 564874 -1644 565494 -1548
rect 579154 597212 579774 598268
rect 579154 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 579774 597212
rect 579154 597088 579774 597156
rect 579154 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 579774 597088
rect 579154 596964 579774 597032
rect 579154 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 579774 596964
rect 579154 596840 579774 596908
rect 579154 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 579774 596840
rect 579154 580350 579774 596784
rect 579154 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 579774 580350
rect 579154 580226 579774 580294
rect 579154 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 579774 580226
rect 579154 580102 579774 580170
rect 579154 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 579774 580102
rect 579154 579978 579774 580046
rect 579154 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 579774 579978
rect 579154 562350 579774 579922
rect 579154 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 579774 562350
rect 579154 562226 579774 562294
rect 579154 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 579774 562226
rect 579154 562102 579774 562170
rect 579154 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 579774 562102
rect 579154 561978 579774 562046
rect 579154 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 579774 561978
rect 579154 544350 579774 561922
rect 579154 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 579774 544350
rect 579154 544226 579774 544294
rect 579154 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 579774 544226
rect 579154 544102 579774 544170
rect 579154 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 579774 544102
rect 579154 543978 579774 544046
rect 579154 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 579774 543978
rect 579154 526350 579774 543922
rect 579154 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 579774 526350
rect 579154 526226 579774 526294
rect 579154 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 579774 526226
rect 579154 526102 579774 526170
rect 579154 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 579774 526102
rect 579154 525978 579774 526046
rect 579154 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 579774 525978
rect 579154 508350 579774 525922
rect 579154 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 579774 508350
rect 579154 508226 579774 508294
rect 579154 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 579774 508226
rect 579154 508102 579774 508170
rect 579154 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 579774 508102
rect 579154 507978 579774 508046
rect 579154 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 579774 507978
rect 579154 490350 579774 507922
rect 579154 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 579774 490350
rect 579154 490226 579774 490294
rect 579154 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 579774 490226
rect 579154 490102 579774 490170
rect 579154 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 579774 490102
rect 579154 489978 579774 490046
rect 579154 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 579774 489978
rect 579154 472350 579774 489922
rect 579154 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 579774 472350
rect 579154 472226 579774 472294
rect 579154 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 579774 472226
rect 579154 472102 579774 472170
rect 579154 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 579774 472102
rect 579154 471978 579774 472046
rect 579154 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 579774 471978
rect 579154 454350 579774 471922
rect 579154 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 579774 454350
rect 579154 454226 579774 454294
rect 579154 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 579774 454226
rect 579154 454102 579774 454170
rect 579154 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 579774 454102
rect 579154 453978 579774 454046
rect 579154 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 579774 453978
rect 579154 436350 579774 453922
rect 579154 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 579774 436350
rect 579154 436226 579774 436294
rect 579154 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 579774 436226
rect 579154 436102 579774 436170
rect 579154 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 579774 436102
rect 579154 435978 579774 436046
rect 579154 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 579774 435978
rect 579154 418350 579774 435922
rect 579154 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 579774 418350
rect 579154 418226 579774 418294
rect 579154 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 579774 418226
rect 579154 418102 579774 418170
rect 579154 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 579774 418102
rect 579154 417978 579774 418046
rect 579154 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 579774 417978
rect 579154 400350 579774 417922
rect 579154 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 579774 400350
rect 579154 400226 579774 400294
rect 579154 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 579774 400226
rect 579154 400102 579774 400170
rect 579154 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 579774 400102
rect 579154 399978 579774 400046
rect 579154 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 579774 399978
rect 579154 382350 579774 399922
rect 579154 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 579774 382350
rect 579154 382226 579774 382294
rect 579154 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 579774 382226
rect 579154 382102 579774 382170
rect 579154 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 579774 382102
rect 579154 381978 579774 382046
rect 579154 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 579774 381978
rect 579154 364350 579774 381922
rect 579154 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 579774 364350
rect 579154 364226 579774 364294
rect 579154 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 579774 364226
rect 579154 364102 579774 364170
rect 579154 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 579774 364102
rect 579154 363978 579774 364046
rect 579154 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 579774 363978
rect 579154 346350 579774 363922
rect 579154 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 579774 346350
rect 579154 346226 579774 346294
rect 579154 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 579774 346226
rect 579154 346102 579774 346170
rect 579154 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 579774 346102
rect 579154 345978 579774 346046
rect 579154 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 579774 345978
rect 579154 328350 579774 345922
rect 579154 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 579774 328350
rect 579154 328226 579774 328294
rect 579154 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 579774 328226
rect 579154 328102 579774 328170
rect 579154 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 579774 328102
rect 579154 327978 579774 328046
rect 579154 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 579774 327978
rect 579154 310350 579774 327922
rect 579154 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 579774 310350
rect 579154 310226 579774 310294
rect 579154 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 579774 310226
rect 579154 310102 579774 310170
rect 579154 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 579774 310102
rect 579154 309978 579774 310046
rect 579154 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 579774 309978
rect 579154 292350 579774 309922
rect 579154 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 579774 292350
rect 579154 292226 579774 292294
rect 579154 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 579774 292226
rect 579154 292102 579774 292170
rect 579154 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 579774 292102
rect 579154 291978 579774 292046
rect 579154 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 579774 291978
rect 579154 274350 579774 291922
rect 579154 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 579774 274350
rect 579154 274226 579774 274294
rect 579154 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 579774 274226
rect 579154 274102 579774 274170
rect 579154 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 579774 274102
rect 579154 273978 579774 274046
rect 579154 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 579774 273978
rect 579154 256350 579774 273922
rect 579154 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 579774 256350
rect 579154 256226 579774 256294
rect 579154 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 579774 256226
rect 579154 256102 579774 256170
rect 579154 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 579774 256102
rect 579154 255978 579774 256046
rect 579154 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 579774 255978
rect 579154 238350 579774 255922
rect 579154 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 579774 238350
rect 579154 238226 579774 238294
rect 579154 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 579774 238226
rect 579154 238102 579774 238170
rect 579154 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 579774 238102
rect 579154 237978 579774 238046
rect 579154 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 579774 237978
rect 579154 220350 579774 237922
rect 579154 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 579774 220350
rect 579154 220226 579774 220294
rect 579154 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 579774 220226
rect 579154 220102 579774 220170
rect 579154 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 579774 220102
rect 579154 219978 579774 220046
rect 579154 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 579774 219978
rect 579154 202350 579774 219922
rect 579154 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 579774 202350
rect 579154 202226 579774 202294
rect 579154 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 579774 202226
rect 579154 202102 579774 202170
rect 579154 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 579774 202102
rect 579154 201978 579774 202046
rect 579154 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 579774 201978
rect 579154 184350 579774 201922
rect 579154 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 579774 184350
rect 579154 184226 579774 184294
rect 579154 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 579774 184226
rect 579154 184102 579774 184170
rect 579154 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 579774 184102
rect 579154 183978 579774 184046
rect 579154 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 579774 183978
rect 579154 166350 579774 183922
rect 579154 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 579774 166350
rect 579154 166226 579774 166294
rect 579154 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 579774 166226
rect 579154 166102 579774 166170
rect 579154 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 579774 166102
rect 579154 165978 579774 166046
rect 579154 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 579774 165978
rect 579154 148350 579774 165922
rect 579154 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 579774 148350
rect 579154 148226 579774 148294
rect 579154 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 579774 148226
rect 579154 148102 579774 148170
rect 579154 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 579774 148102
rect 579154 147978 579774 148046
rect 579154 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 579774 147978
rect 579154 130350 579774 147922
rect 579154 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 579774 130350
rect 579154 130226 579774 130294
rect 579154 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 579774 130226
rect 579154 130102 579774 130170
rect 579154 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 579774 130102
rect 579154 129978 579774 130046
rect 579154 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 579774 129978
rect 579154 112350 579774 129922
rect 579154 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 579774 112350
rect 579154 112226 579774 112294
rect 579154 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 579774 112226
rect 579154 112102 579774 112170
rect 579154 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 579774 112102
rect 579154 111978 579774 112046
rect 579154 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 579774 111978
rect 579154 94350 579774 111922
rect 579154 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 579774 94350
rect 579154 94226 579774 94294
rect 579154 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 579774 94226
rect 579154 94102 579774 94170
rect 579154 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 579774 94102
rect 579154 93978 579774 94046
rect 579154 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 579774 93978
rect 579154 76350 579774 93922
rect 579154 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 579774 76350
rect 579154 76226 579774 76294
rect 579154 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 579774 76226
rect 579154 76102 579774 76170
rect 579154 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 579774 76102
rect 579154 75978 579774 76046
rect 579154 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 579774 75978
rect 579154 58350 579774 75922
rect 579154 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 579774 58350
rect 579154 58226 579774 58294
rect 579154 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 579774 58226
rect 579154 58102 579774 58170
rect 579154 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 579774 58102
rect 579154 57978 579774 58046
rect 579154 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 579774 57978
rect 579154 40350 579774 57922
rect 579154 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 579774 40350
rect 579154 40226 579774 40294
rect 579154 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 579774 40226
rect 579154 40102 579774 40170
rect 579154 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 579774 40102
rect 579154 39978 579774 40046
rect 579154 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 579774 39978
rect 579154 22350 579774 39922
rect 579154 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 579774 22350
rect 579154 22226 579774 22294
rect 579154 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 579774 22226
rect 579154 22102 579774 22170
rect 579154 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 579774 22102
rect 579154 21978 579774 22046
rect 579154 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 579774 21978
rect 579154 4350 579774 21922
rect 579154 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 579774 4350
rect 579154 4226 579774 4294
rect 579154 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 579774 4226
rect 579154 4102 579774 4170
rect 579154 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 579774 4102
rect 579154 3978 579774 4046
rect 579154 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 579774 3978
rect 579154 -160 579774 3922
rect 579154 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 579774 -160
rect 579154 -284 579774 -216
rect 579154 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 579774 -284
rect 579154 -408 579774 -340
rect 579154 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 579774 -408
rect 579154 -532 579774 -464
rect 579154 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 579774 -532
rect 579154 -1644 579774 -588
rect 582874 598172 583494 598268
rect 582874 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 583494 598172
rect 582874 598048 583494 598116
rect 582874 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 583494 598048
rect 582874 597924 583494 597992
rect 582874 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 583494 597924
rect 582874 597800 583494 597868
rect 582874 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 583494 597800
rect 582874 586350 583494 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 582874 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 583494 586350
rect 582874 586226 583494 586294
rect 582874 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 583494 586226
rect 582874 586102 583494 586170
rect 582874 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 583494 586102
rect 582874 585978 583494 586046
rect 582874 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 583494 585978
rect 582874 568350 583494 585922
rect 582874 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 583494 568350
rect 582874 568226 583494 568294
rect 582874 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 583494 568226
rect 582874 568102 583494 568170
rect 582874 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 583494 568102
rect 582874 567978 583494 568046
rect 582874 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 583494 567978
rect 582874 550350 583494 567922
rect 582874 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 583494 550350
rect 582874 550226 583494 550294
rect 582874 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 583494 550226
rect 582874 550102 583494 550170
rect 582874 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 583494 550102
rect 582874 549978 583494 550046
rect 582874 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 583494 549978
rect 582874 532350 583494 549922
rect 582874 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 583494 532350
rect 582874 532226 583494 532294
rect 582874 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 583494 532226
rect 582874 532102 583494 532170
rect 582874 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 583494 532102
rect 582874 531978 583494 532046
rect 582874 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 583494 531978
rect 582874 514350 583494 531922
rect 582874 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 583494 514350
rect 582874 514226 583494 514294
rect 582874 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 583494 514226
rect 582874 514102 583494 514170
rect 582874 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 583494 514102
rect 582874 513978 583494 514046
rect 582874 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 583494 513978
rect 582874 496350 583494 513922
rect 582874 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 583494 496350
rect 582874 496226 583494 496294
rect 582874 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 583494 496226
rect 582874 496102 583494 496170
rect 582874 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 583494 496102
rect 582874 495978 583494 496046
rect 582874 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 583494 495978
rect 582874 478350 583494 495922
rect 582874 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 583494 478350
rect 582874 478226 583494 478294
rect 582874 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 583494 478226
rect 582874 478102 583494 478170
rect 582874 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 583494 478102
rect 582874 477978 583494 478046
rect 582874 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 583494 477978
rect 582874 460350 583494 477922
rect 582874 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 583494 460350
rect 582874 460226 583494 460294
rect 582874 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 583494 460226
rect 582874 460102 583494 460170
rect 582874 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 583494 460102
rect 582874 459978 583494 460046
rect 582874 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 583494 459978
rect 582874 442350 583494 459922
rect 582874 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 583494 442350
rect 582874 442226 583494 442294
rect 582874 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 583494 442226
rect 582874 442102 583494 442170
rect 582874 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 583494 442102
rect 582874 441978 583494 442046
rect 582874 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 583494 441978
rect 582874 424350 583494 441922
rect 582874 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 583494 424350
rect 582874 424226 583494 424294
rect 582874 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 583494 424226
rect 582874 424102 583494 424170
rect 582874 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 583494 424102
rect 582874 423978 583494 424046
rect 582874 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 583494 423978
rect 582874 406350 583494 423922
rect 582874 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 583494 406350
rect 582874 406226 583494 406294
rect 582874 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 583494 406226
rect 582874 406102 583494 406170
rect 582874 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 583494 406102
rect 582874 405978 583494 406046
rect 582874 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 583494 405978
rect 582874 388350 583494 405922
rect 582874 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 583494 388350
rect 582874 388226 583494 388294
rect 582874 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 583494 388226
rect 582874 388102 583494 388170
rect 582874 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 583494 388102
rect 582874 387978 583494 388046
rect 582874 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 583494 387978
rect 582874 370350 583494 387922
rect 582874 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 583494 370350
rect 582874 370226 583494 370294
rect 582874 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 583494 370226
rect 582874 370102 583494 370170
rect 582874 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 583494 370102
rect 582874 369978 583494 370046
rect 582874 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 583494 369978
rect 582874 352350 583494 369922
rect 582874 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 583494 352350
rect 582874 352226 583494 352294
rect 582874 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 583494 352226
rect 582874 352102 583494 352170
rect 582874 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 583494 352102
rect 582874 351978 583494 352046
rect 582874 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 583494 351978
rect 582874 334350 583494 351922
rect 582874 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 583494 334350
rect 582874 334226 583494 334294
rect 582874 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 583494 334226
rect 582874 334102 583494 334170
rect 582874 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 583494 334102
rect 582874 333978 583494 334046
rect 582874 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 583494 333978
rect 582874 316350 583494 333922
rect 582874 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 583494 316350
rect 582874 316226 583494 316294
rect 582874 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 583494 316226
rect 582874 316102 583494 316170
rect 582874 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 583494 316102
rect 582874 315978 583494 316046
rect 582874 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 583494 315978
rect 582874 298350 583494 315922
rect 582874 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 583494 298350
rect 582874 298226 583494 298294
rect 582874 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 583494 298226
rect 582874 298102 583494 298170
rect 582874 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 583494 298102
rect 582874 297978 583494 298046
rect 582874 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 583494 297978
rect 582874 280350 583494 297922
rect 582874 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 583494 280350
rect 582874 280226 583494 280294
rect 582874 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 583494 280226
rect 582874 280102 583494 280170
rect 582874 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 583494 280102
rect 582874 279978 583494 280046
rect 582874 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 583494 279978
rect 582874 262350 583494 279922
rect 582874 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 583494 262350
rect 582874 262226 583494 262294
rect 582874 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 583494 262226
rect 582874 262102 583494 262170
rect 582874 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 583494 262102
rect 582874 261978 583494 262046
rect 582874 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 583494 261978
rect 582874 244350 583494 261922
rect 582874 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 583494 244350
rect 582874 244226 583494 244294
rect 582874 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 583494 244226
rect 582874 244102 583494 244170
rect 582874 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 583494 244102
rect 582874 243978 583494 244046
rect 582874 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 583494 243978
rect 582874 226350 583494 243922
rect 582874 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 583494 226350
rect 582874 226226 583494 226294
rect 582874 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 583494 226226
rect 582874 226102 583494 226170
rect 582874 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 583494 226102
rect 582874 225978 583494 226046
rect 582874 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 583494 225978
rect 582874 208350 583494 225922
rect 582874 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 583494 208350
rect 582874 208226 583494 208294
rect 582874 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 583494 208226
rect 582874 208102 583494 208170
rect 582874 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 583494 208102
rect 582874 207978 583494 208046
rect 582874 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 583494 207978
rect 582874 190350 583494 207922
rect 582874 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 583494 190350
rect 582874 190226 583494 190294
rect 582874 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 583494 190226
rect 582874 190102 583494 190170
rect 582874 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 583494 190102
rect 582874 189978 583494 190046
rect 582874 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 583494 189978
rect 582874 172350 583494 189922
rect 582874 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 583494 172350
rect 582874 172226 583494 172294
rect 582874 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 583494 172226
rect 582874 172102 583494 172170
rect 582874 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 583494 172102
rect 582874 171978 583494 172046
rect 582874 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 583494 171978
rect 582874 154350 583494 171922
rect 582874 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 583494 154350
rect 582874 154226 583494 154294
rect 582874 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 583494 154226
rect 582874 154102 583494 154170
rect 582874 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 583494 154102
rect 582874 153978 583494 154046
rect 582874 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 583494 153978
rect 582874 136350 583494 153922
rect 582874 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 583494 136350
rect 582874 136226 583494 136294
rect 582874 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 583494 136226
rect 582874 136102 583494 136170
rect 582874 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 583494 136102
rect 582874 135978 583494 136046
rect 582874 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 583494 135978
rect 582874 118350 583494 135922
rect 582874 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 583494 118350
rect 582874 118226 583494 118294
rect 582874 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 583494 118226
rect 582874 118102 583494 118170
rect 582874 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 583494 118102
rect 582874 117978 583494 118046
rect 582874 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 583494 117978
rect 582874 100350 583494 117922
rect 582874 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 583494 100350
rect 582874 100226 583494 100294
rect 582874 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 583494 100226
rect 582874 100102 583494 100170
rect 582874 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 583494 100102
rect 582874 99978 583494 100046
rect 582874 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 583494 99978
rect 582874 82350 583494 99922
rect 582874 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 583494 82350
rect 582874 82226 583494 82294
rect 582874 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 583494 82226
rect 582874 82102 583494 82170
rect 582874 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 583494 82102
rect 582874 81978 583494 82046
rect 582874 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 583494 81978
rect 582874 64350 583494 81922
rect 582874 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 583494 64350
rect 582874 64226 583494 64294
rect 582874 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 583494 64226
rect 582874 64102 583494 64170
rect 582874 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 583494 64102
rect 582874 63978 583494 64046
rect 582874 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 583494 63978
rect 582874 46350 583494 63922
rect 582874 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 583494 46350
rect 582874 46226 583494 46294
rect 582874 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 583494 46226
rect 582874 46102 583494 46170
rect 582874 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 583494 46102
rect 582874 45978 583494 46046
rect 582874 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 583494 45978
rect 582874 28350 583494 45922
rect 582874 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 583494 28350
rect 582874 28226 583494 28294
rect 582874 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 583494 28226
rect 582874 28102 583494 28170
rect 582874 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 583494 28102
rect 582874 27978 583494 28046
rect 582874 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 583494 27978
rect 582874 10350 583494 27922
rect 582874 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 583494 10350
rect 582874 10226 583494 10294
rect 582874 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 583494 10226
rect 582874 10102 583494 10170
rect 582874 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 583494 10102
rect 582874 9978 583494 10046
rect 582874 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 583494 9978
rect 582874 -1120 583494 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 582874 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 583494 -1120
rect 582874 -1244 583494 -1176
rect 582874 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 583494 -1244
rect 582874 -1368 583494 -1300
rect 582874 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 583494 -1368
rect 582874 -1492 583494 -1424
rect 582874 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 583494 -1492
rect 582874 -1644 583494 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 3250 597156 3306 597212
rect 3374 597156 3430 597212
rect 3498 597156 3554 597212
rect 3622 597156 3678 597212
rect 3250 597032 3306 597088
rect 3374 597032 3430 597088
rect 3498 597032 3554 597088
rect 3622 597032 3678 597088
rect 3250 596908 3306 596964
rect 3374 596908 3430 596964
rect 3498 596908 3554 596964
rect 3622 596908 3678 596964
rect 3250 596784 3306 596840
rect 3374 596784 3430 596840
rect 3498 596784 3554 596840
rect 3622 596784 3678 596840
rect 3250 580294 3306 580350
rect 3374 580294 3430 580350
rect 3498 580294 3554 580350
rect 3622 580294 3678 580350
rect 3250 580170 3306 580226
rect 3374 580170 3430 580226
rect 3498 580170 3554 580226
rect 3622 580170 3678 580226
rect 3250 580046 3306 580102
rect 3374 580046 3430 580102
rect 3498 580046 3554 580102
rect 3622 580046 3678 580102
rect 3250 579922 3306 579978
rect 3374 579922 3430 579978
rect 3498 579922 3554 579978
rect 3622 579922 3678 579978
rect 3250 562294 3306 562350
rect 3374 562294 3430 562350
rect 3498 562294 3554 562350
rect 3622 562294 3678 562350
rect 3250 562170 3306 562226
rect 3374 562170 3430 562226
rect 3498 562170 3554 562226
rect 3622 562170 3678 562226
rect 3250 562046 3306 562102
rect 3374 562046 3430 562102
rect 3498 562046 3554 562102
rect 3622 562046 3678 562102
rect 3250 561922 3306 561978
rect 3374 561922 3430 561978
rect 3498 561922 3554 561978
rect 3622 561922 3678 561978
rect 3250 544294 3306 544350
rect 3374 544294 3430 544350
rect 3498 544294 3554 544350
rect 3622 544294 3678 544350
rect 3250 544170 3306 544226
rect 3374 544170 3430 544226
rect 3498 544170 3554 544226
rect 3622 544170 3678 544226
rect 3250 544046 3306 544102
rect 3374 544046 3430 544102
rect 3498 544046 3554 544102
rect 3622 544046 3678 544102
rect 3250 543922 3306 543978
rect 3374 543922 3430 543978
rect 3498 543922 3554 543978
rect 3622 543922 3678 543978
rect 3250 526294 3306 526350
rect 3374 526294 3430 526350
rect 3498 526294 3554 526350
rect 3622 526294 3678 526350
rect 3250 526170 3306 526226
rect 3374 526170 3430 526226
rect 3498 526170 3554 526226
rect 3622 526170 3678 526226
rect 3250 526046 3306 526102
rect 3374 526046 3430 526102
rect 3498 526046 3554 526102
rect 3622 526046 3678 526102
rect 3250 525922 3306 525978
rect 3374 525922 3430 525978
rect 3498 525922 3554 525978
rect 3622 525922 3678 525978
rect 3250 508294 3306 508350
rect 3374 508294 3430 508350
rect 3498 508294 3554 508350
rect 3622 508294 3678 508350
rect 3250 508170 3306 508226
rect 3374 508170 3430 508226
rect 3498 508170 3554 508226
rect 3622 508170 3678 508226
rect 3250 508046 3306 508102
rect 3374 508046 3430 508102
rect 3498 508046 3554 508102
rect 3622 508046 3678 508102
rect 3250 507922 3306 507978
rect 3374 507922 3430 507978
rect 3498 507922 3554 507978
rect 3622 507922 3678 507978
rect 3250 490294 3306 490350
rect 3374 490294 3430 490350
rect 3498 490294 3554 490350
rect 3622 490294 3678 490350
rect 3250 490170 3306 490226
rect 3374 490170 3430 490226
rect 3498 490170 3554 490226
rect 3622 490170 3678 490226
rect 3250 490046 3306 490102
rect 3374 490046 3430 490102
rect 3498 490046 3554 490102
rect 3622 490046 3678 490102
rect 3250 489922 3306 489978
rect 3374 489922 3430 489978
rect 3498 489922 3554 489978
rect 3622 489922 3678 489978
rect 3250 472294 3306 472350
rect 3374 472294 3430 472350
rect 3498 472294 3554 472350
rect 3622 472294 3678 472350
rect 3250 472170 3306 472226
rect 3374 472170 3430 472226
rect 3498 472170 3554 472226
rect 3622 472170 3678 472226
rect 3250 472046 3306 472102
rect 3374 472046 3430 472102
rect 3498 472046 3554 472102
rect 3622 472046 3678 472102
rect 3250 471922 3306 471978
rect 3374 471922 3430 471978
rect 3498 471922 3554 471978
rect 3622 471922 3678 471978
rect 3250 454294 3306 454350
rect 3374 454294 3430 454350
rect 3498 454294 3554 454350
rect 3622 454294 3678 454350
rect 3250 454170 3306 454226
rect 3374 454170 3430 454226
rect 3498 454170 3554 454226
rect 3622 454170 3678 454226
rect 3250 454046 3306 454102
rect 3374 454046 3430 454102
rect 3498 454046 3554 454102
rect 3622 454046 3678 454102
rect 3250 453922 3306 453978
rect 3374 453922 3430 453978
rect 3498 453922 3554 453978
rect 3622 453922 3678 453978
rect 3250 436294 3306 436350
rect 3374 436294 3430 436350
rect 3498 436294 3554 436350
rect 3622 436294 3678 436350
rect 3250 436170 3306 436226
rect 3374 436170 3430 436226
rect 3498 436170 3554 436226
rect 3622 436170 3678 436226
rect 3250 436046 3306 436102
rect 3374 436046 3430 436102
rect 3498 436046 3554 436102
rect 3622 436046 3678 436102
rect 3250 435922 3306 435978
rect 3374 435922 3430 435978
rect 3498 435922 3554 435978
rect 3622 435922 3678 435978
rect 3250 418294 3306 418350
rect 3374 418294 3430 418350
rect 3498 418294 3554 418350
rect 3622 418294 3678 418350
rect 3250 418170 3306 418226
rect 3374 418170 3430 418226
rect 3498 418170 3554 418226
rect 3622 418170 3678 418226
rect 3250 418046 3306 418102
rect 3374 418046 3430 418102
rect 3498 418046 3554 418102
rect 3622 418046 3678 418102
rect 3250 417922 3306 417978
rect 3374 417922 3430 417978
rect 3498 417922 3554 417978
rect 3622 417922 3678 417978
rect 3250 400294 3306 400350
rect 3374 400294 3430 400350
rect 3498 400294 3554 400350
rect 3622 400294 3678 400350
rect 3250 400170 3306 400226
rect 3374 400170 3430 400226
rect 3498 400170 3554 400226
rect 3622 400170 3678 400226
rect 3250 400046 3306 400102
rect 3374 400046 3430 400102
rect 3498 400046 3554 400102
rect 3622 400046 3678 400102
rect 3250 399922 3306 399978
rect 3374 399922 3430 399978
rect 3498 399922 3554 399978
rect 3622 399922 3678 399978
rect 3250 382294 3306 382350
rect 3374 382294 3430 382350
rect 3498 382294 3554 382350
rect 3622 382294 3678 382350
rect 3250 382170 3306 382226
rect 3374 382170 3430 382226
rect 3498 382170 3554 382226
rect 3622 382170 3678 382226
rect 3250 382046 3306 382102
rect 3374 382046 3430 382102
rect 3498 382046 3554 382102
rect 3622 382046 3678 382102
rect 3250 381922 3306 381978
rect 3374 381922 3430 381978
rect 3498 381922 3554 381978
rect 3622 381922 3678 381978
rect 3250 364294 3306 364350
rect 3374 364294 3430 364350
rect 3498 364294 3554 364350
rect 3622 364294 3678 364350
rect 3250 364170 3306 364226
rect 3374 364170 3430 364226
rect 3498 364170 3554 364226
rect 3622 364170 3678 364226
rect 3250 364046 3306 364102
rect 3374 364046 3430 364102
rect 3498 364046 3554 364102
rect 3622 364046 3678 364102
rect 3250 363922 3306 363978
rect 3374 363922 3430 363978
rect 3498 363922 3554 363978
rect 3622 363922 3678 363978
rect 3250 346294 3306 346350
rect 3374 346294 3430 346350
rect 3498 346294 3554 346350
rect 3622 346294 3678 346350
rect 3250 346170 3306 346226
rect 3374 346170 3430 346226
rect 3498 346170 3554 346226
rect 3622 346170 3678 346226
rect 3250 346046 3306 346102
rect 3374 346046 3430 346102
rect 3498 346046 3554 346102
rect 3622 346046 3678 346102
rect 3250 345922 3306 345978
rect 3374 345922 3430 345978
rect 3498 345922 3554 345978
rect 3622 345922 3678 345978
rect 3250 328294 3306 328350
rect 3374 328294 3430 328350
rect 3498 328294 3554 328350
rect 3622 328294 3678 328350
rect 3250 328170 3306 328226
rect 3374 328170 3430 328226
rect 3498 328170 3554 328226
rect 3622 328170 3678 328226
rect 3250 328046 3306 328102
rect 3374 328046 3430 328102
rect 3498 328046 3554 328102
rect 3622 328046 3678 328102
rect 3250 327922 3306 327978
rect 3374 327922 3430 327978
rect 3498 327922 3554 327978
rect 3622 327922 3678 327978
rect 3250 310294 3306 310350
rect 3374 310294 3430 310350
rect 3498 310294 3554 310350
rect 3622 310294 3678 310350
rect 3250 310170 3306 310226
rect 3374 310170 3430 310226
rect 3498 310170 3554 310226
rect 3622 310170 3678 310226
rect 3250 310046 3306 310102
rect 3374 310046 3430 310102
rect 3498 310046 3554 310102
rect 3622 310046 3678 310102
rect 3250 309922 3306 309978
rect 3374 309922 3430 309978
rect 3498 309922 3554 309978
rect 3622 309922 3678 309978
rect 3250 292294 3306 292350
rect 3374 292294 3430 292350
rect 3498 292294 3554 292350
rect 3622 292294 3678 292350
rect 3250 292170 3306 292226
rect 3374 292170 3430 292226
rect 3498 292170 3554 292226
rect 3622 292170 3678 292226
rect 3250 292046 3306 292102
rect 3374 292046 3430 292102
rect 3498 292046 3554 292102
rect 3622 292046 3678 292102
rect 3250 291922 3306 291978
rect 3374 291922 3430 291978
rect 3498 291922 3554 291978
rect 3622 291922 3678 291978
rect 3250 274294 3306 274350
rect 3374 274294 3430 274350
rect 3498 274294 3554 274350
rect 3622 274294 3678 274350
rect 3250 274170 3306 274226
rect 3374 274170 3430 274226
rect 3498 274170 3554 274226
rect 3622 274170 3678 274226
rect 3250 274046 3306 274102
rect 3374 274046 3430 274102
rect 3498 274046 3554 274102
rect 3622 274046 3678 274102
rect 3250 273922 3306 273978
rect 3374 273922 3430 273978
rect 3498 273922 3554 273978
rect 3622 273922 3678 273978
rect 3250 256294 3306 256350
rect 3374 256294 3430 256350
rect 3498 256294 3554 256350
rect 3622 256294 3678 256350
rect 3250 256170 3306 256226
rect 3374 256170 3430 256226
rect 3498 256170 3554 256226
rect 3622 256170 3678 256226
rect 3250 256046 3306 256102
rect 3374 256046 3430 256102
rect 3498 256046 3554 256102
rect 3622 256046 3678 256102
rect 3250 255922 3306 255978
rect 3374 255922 3430 255978
rect 3498 255922 3554 255978
rect 3622 255922 3678 255978
rect 3250 238294 3306 238350
rect 3374 238294 3430 238350
rect 3498 238294 3554 238350
rect 3622 238294 3678 238350
rect 3250 238170 3306 238226
rect 3374 238170 3430 238226
rect 3498 238170 3554 238226
rect 3622 238170 3678 238226
rect 3250 238046 3306 238102
rect 3374 238046 3430 238102
rect 3498 238046 3554 238102
rect 3622 238046 3678 238102
rect 3250 237922 3306 237978
rect 3374 237922 3430 237978
rect 3498 237922 3554 237978
rect 3622 237922 3678 237978
rect 3250 220294 3306 220350
rect 3374 220294 3430 220350
rect 3498 220294 3554 220350
rect 3622 220294 3678 220350
rect 3250 220170 3306 220226
rect 3374 220170 3430 220226
rect 3498 220170 3554 220226
rect 3622 220170 3678 220226
rect 3250 220046 3306 220102
rect 3374 220046 3430 220102
rect 3498 220046 3554 220102
rect 3622 220046 3678 220102
rect 3250 219922 3306 219978
rect 3374 219922 3430 219978
rect 3498 219922 3554 219978
rect 3622 219922 3678 219978
rect 3250 202294 3306 202350
rect 3374 202294 3430 202350
rect 3498 202294 3554 202350
rect 3622 202294 3678 202350
rect 3250 202170 3306 202226
rect 3374 202170 3430 202226
rect 3498 202170 3554 202226
rect 3622 202170 3678 202226
rect 3250 202046 3306 202102
rect 3374 202046 3430 202102
rect 3498 202046 3554 202102
rect 3622 202046 3678 202102
rect 3250 201922 3306 201978
rect 3374 201922 3430 201978
rect 3498 201922 3554 201978
rect 3622 201922 3678 201978
rect 3250 184294 3306 184350
rect 3374 184294 3430 184350
rect 3498 184294 3554 184350
rect 3622 184294 3678 184350
rect 3250 184170 3306 184226
rect 3374 184170 3430 184226
rect 3498 184170 3554 184226
rect 3622 184170 3678 184226
rect 3250 184046 3306 184102
rect 3374 184046 3430 184102
rect 3498 184046 3554 184102
rect 3622 184046 3678 184102
rect 3250 183922 3306 183978
rect 3374 183922 3430 183978
rect 3498 183922 3554 183978
rect 3622 183922 3678 183978
rect 3250 166294 3306 166350
rect 3374 166294 3430 166350
rect 3498 166294 3554 166350
rect 3622 166294 3678 166350
rect 3250 166170 3306 166226
rect 3374 166170 3430 166226
rect 3498 166170 3554 166226
rect 3622 166170 3678 166226
rect 3250 166046 3306 166102
rect 3374 166046 3430 166102
rect 3498 166046 3554 166102
rect 3622 166046 3678 166102
rect 3250 165922 3306 165978
rect 3374 165922 3430 165978
rect 3498 165922 3554 165978
rect 3622 165922 3678 165978
rect 3250 148294 3306 148350
rect 3374 148294 3430 148350
rect 3498 148294 3554 148350
rect 3622 148294 3678 148350
rect 3250 148170 3306 148226
rect 3374 148170 3430 148226
rect 3498 148170 3554 148226
rect 3622 148170 3678 148226
rect 3250 148046 3306 148102
rect 3374 148046 3430 148102
rect 3498 148046 3554 148102
rect 3622 148046 3678 148102
rect 3250 147922 3306 147978
rect 3374 147922 3430 147978
rect 3498 147922 3554 147978
rect 3622 147922 3678 147978
rect 3250 130294 3306 130350
rect 3374 130294 3430 130350
rect 3498 130294 3554 130350
rect 3622 130294 3678 130350
rect 3250 130170 3306 130226
rect 3374 130170 3430 130226
rect 3498 130170 3554 130226
rect 3622 130170 3678 130226
rect 3250 130046 3306 130102
rect 3374 130046 3430 130102
rect 3498 130046 3554 130102
rect 3622 130046 3678 130102
rect 3250 129922 3306 129978
rect 3374 129922 3430 129978
rect 3498 129922 3554 129978
rect 3622 129922 3678 129978
rect 3250 112294 3306 112350
rect 3374 112294 3430 112350
rect 3498 112294 3554 112350
rect 3622 112294 3678 112350
rect 3250 112170 3306 112226
rect 3374 112170 3430 112226
rect 3498 112170 3554 112226
rect 3622 112170 3678 112226
rect 3250 112046 3306 112102
rect 3374 112046 3430 112102
rect 3498 112046 3554 112102
rect 3622 112046 3678 112102
rect 3250 111922 3306 111978
rect 3374 111922 3430 111978
rect 3498 111922 3554 111978
rect 3622 111922 3678 111978
rect 3250 94294 3306 94350
rect 3374 94294 3430 94350
rect 3498 94294 3554 94350
rect 3622 94294 3678 94350
rect 3250 94170 3306 94226
rect 3374 94170 3430 94226
rect 3498 94170 3554 94226
rect 3622 94170 3678 94226
rect 3250 94046 3306 94102
rect 3374 94046 3430 94102
rect 3498 94046 3554 94102
rect 3622 94046 3678 94102
rect 3250 93922 3306 93978
rect 3374 93922 3430 93978
rect 3498 93922 3554 93978
rect 3622 93922 3678 93978
rect 3250 76294 3306 76350
rect 3374 76294 3430 76350
rect 3498 76294 3554 76350
rect 3622 76294 3678 76350
rect 3250 76170 3306 76226
rect 3374 76170 3430 76226
rect 3498 76170 3554 76226
rect 3622 76170 3678 76226
rect 3250 76046 3306 76102
rect 3374 76046 3430 76102
rect 3498 76046 3554 76102
rect 3622 76046 3678 76102
rect 3250 75922 3306 75978
rect 3374 75922 3430 75978
rect 3498 75922 3554 75978
rect 3622 75922 3678 75978
rect 3250 58294 3306 58350
rect 3374 58294 3430 58350
rect 3498 58294 3554 58350
rect 3622 58294 3678 58350
rect 3250 58170 3306 58226
rect 3374 58170 3430 58226
rect 3498 58170 3554 58226
rect 3622 58170 3678 58226
rect 3250 58046 3306 58102
rect 3374 58046 3430 58102
rect 3498 58046 3554 58102
rect 3622 58046 3678 58102
rect 3250 57922 3306 57978
rect 3374 57922 3430 57978
rect 3498 57922 3554 57978
rect 3622 57922 3678 57978
rect 3250 40294 3306 40350
rect 3374 40294 3430 40350
rect 3498 40294 3554 40350
rect 3622 40294 3678 40350
rect 3250 40170 3306 40226
rect 3374 40170 3430 40226
rect 3498 40170 3554 40226
rect 3622 40170 3678 40226
rect 3250 40046 3306 40102
rect 3374 40046 3430 40102
rect 3498 40046 3554 40102
rect 3622 40046 3678 40102
rect 3250 39922 3306 39978
rect 3374 39922 3430 39978
rect 3498 39922 3554 39978
rect 3622 39922 3678 39978
rect 3250 22294 3306 22350
rect 3374 22294 3430 22350
rect 3498 22294 3554 22350
rect 3622 22294 3678 22350
rect 3250 22170 3306 22226
rect 3374 22170 3430 22226
rect 3498 22170 3554 22226
rect 3622 22170 3678 22226
rect 3250 22046 3306 22102
rect 3374 22046 3430 22102
rect 3498 22046 3554 22102
rect 3622 22046 3678 22102
rect 3250 21922 3306 21978
rect 3374 21922 3430 21978
rect 3498 21922 3554 21978
rect 3622 21922 3678 21978
rect 3250 4294 3306 4350
rect 3374 4294 3430 4350
rect 3498 4294 3554 4350
rect 3622 4294 3678 4350
rect 3250 4170 3306 4226
rect 3374 4170 3430 4226
rect 3498 4170 3554 4226
rect 3622 4170 3678 4226
rect 3250 4046 3306 4102
rect 3374 4046 3430 4102
rect 3498 4046 3554 4102
rect 3622 4046 3678 4102
rect 3250 3922 3306 3978
rect 3374 3922 3430 3978
rect 3498 3922 3554 3978
rect 3622 3922 3678 3978
rect 3250 -216 3306 -160
rect 3374 -216 3430 -160
rect 3498 -216 3554 -160
rect 3622 -216 3678 -160
rect 3250 -340 3306 -284
rect 3374 -340 3430 -284
rect 3498 -340 3554 -284
rect 3622 -340 3678 -284
rect 3250 -464 3306 -408
rect 3374 -464 3430 -408
rect 3498 -464 3554 -408
rect 3622 -464 3678 -408
rect 3250 -588 3306 -532
rect 3374 -588 3430 -532
rect 3498 -588 3554 -532
rect 3622 -588 3678 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 6970 598116 7026 598172
rect 7094 598116 7150 598172
rect 7218 598116 7274 598172
rect 7342 598116 7398 598172
rect 6970 597992 7026 598048
rect 7094 597992 7150 598048
rect 7218 597992 7274 598048
rect 7342 597992 7398 598048
rect 6970 597868 7026 597924
rect 7094 597868 7150 597924
rect 7218 597868 7274 597924
rect 7342 597868 7398 597924
rect 6970 597744 7026 597800
rect 7094 597744 7150 597800
rect 7218 597744 7274 597800
rect 7342 597744 7398 597800
rect 6970 586294 7026 586350
rect 7094 586294 7150 586350
rect 7218 586294 7274 586350
rect 7342 586294 7398 586350
rect 6970 586170 7026 586226
rect 7094 586170 7150 586226
rect 7218 586170 7274 586226
rect 7342 586170 7398 586226
rect 6970 586046 7026 586102
rect 7094 586046 7150 586102
rect 7218 586046 7274 586102
rect 7342 586046 7398 586102
rect 6970 585922 7026 585978
rect 7094 585922 7150 585978
rect 7218 585922 7274 585978
rect 7342 585922 7398 585978
rect 6970 568294 7026 568350
rect 7094 568294 7150 568350
rect 7218 568294 7274 568350
rect 7342 568294 7398 568350
rect 6970 568170 7026 568226
rect 7094 568170 7150 568226
rect 7218 568170 7274 568226
rect 7342 568170 7398 568226
rect 6970 568046 7026 568102
rect 7094 568046 7150 568102
rect 7218 568046 7274 568102
rect 7342 568046 7398 568102
rect 6970 567922 7026 567978
rect 7094 567922 7150 567978
rect 7218 567922 7274 567978
rect 7342 567922 7398 567978
rect 6970 550294 7026 550350
rect 7094 550294 7150 550350
rect 7218 550294 7274 550350
rect 7342 550294 7398 550350
rect 6970 550170 7026 550226
rect 7094 550170 7150 550226
rect 7218 550170 7274 550226
rect 7342 550170 7398 550226
rect 6970 550046 7026 550102
rect 7094 550046 7150 550102
rect 7218 550046 7274 550102
rect 7342 550046 7398 550102
rect 6970 549922 7026 549978
rect 7094 549922 7150 549978
rect 7218 549922 7274 549978
rect 7342 549922 7398 549978
rect 6970 532294 7026 532350
rect 7094 532294 7150 532350
rect 7218 532294 7274 532350
rect 7342 532294 7398 532350
rect 6970 532170 7026 532226
rect 7094 532170 7150 532226
rect 7218 532170 7274 532226
rect 7342 532170 7398 532226
rect 6970 532046 7026 532102
rect 7094 532046 7150 532102
rect 7218 532046 7274 532102
rect 7342 532046 7398 532102
rect 6970 531922 7026 531978
rect 7094 531922 7150 531978
rect 7218 531922 7274 531978
rect 7342 531922 7398 531978
rect 21250 597156 21306 597212
rect 21374 597156 21430 597212
rect 21498 597156 21554 597212
rect 21622 597156 21678 597212
rect 21250 597032 21306 597088
rect 21374 597032 21430 597088
rect 21498 597032 21554 597088
rect 21622 597032 21678 597088
rect 21250 596908 21306 596964
rect 21374 596908 21430 596964
rect 21498 596908 21554 596964
rect 21622 596908 21678 596964
rect 21250 596784 21306 596840
rect 21374 596784 21430 596840
rect 21498 596784 21554 596840
rect 21622 596784 21678 596840
rect 21250 580294 21306 580350
rect 21374 580294 21430 580350
rect 21498 580294 21554 580350
rect 21622 580294 21678 580350
rect 21250 580170 21306 580226
rect 21374 580170 21430 580226
rect 21498 580170 21554 580226
rect 21622 580170 21678 580226
rect 21250 580046 21306 580102
rect 21374 580046 21430 580102
rect 21498 580046 21554 580102
rect 21622 580046 21678 580102
rect 21250 579922 21306 579978
rect 21374 579922 21430 579978
rect 21498 579922 21554 579978
rect 21622 579922 21678 579978
rect 21250 562294 21306 562350
rect 21374 562294 21430 562350
rect 21498 562294 21554 562350
rect 21622 562294 21678 562350
rect 21250 562170 21306 562226
rect 21374 562170 21430 562226
rect 21498 562170 21554 562226
rect 21622 562170 21678 562226
rect 21250 562046 21306 562102
rect 21374 562046 21430 562102
rect 21498 562046 21554 562102
rect 21622 562046 21678 562102
rect 21250 561922 21306 561978
rect 21374 561922 21430 561978
rect 21498 561922 21554 561978
rect 21622 561922 21678 561978
rect 21250 544294 21306 544350
rect 21374 544294 21430 544350
rect 21498 544294 21554 544350
rect 21622 544294 21678 544350
rect 21250 544170 21306 544226
rect 21374 544170 21430 544226
rect 21498 544170 21554 544226
rect 21622 544170 21678 544226
rect 21250 544046 21306 544102
rect 21374 544046 21430 544102
rect 21498 544046 21554 544102
rect 21622 544046 21678 544102
rect 21250 543922 21306 543978
rect 21374 543922 21430 543978
rect 21498 543922 21554 543978
rect 21622 543922 21678 543978
rect 21250 526294 21306 526350
rect 21374 526294 21430 526350
rect 21498 526294 21554 526350
rect 21622 526294 21678 526350
rect 21250 526170 21306 526226
rect 21374 526170 21430 526226
rect 21498 526170 21554 526226
rect 21622 526170 21678 526226
rect 21250 526046 21306 526102
rect 21374 526046 21430 526102
rect 21498 526046 21554 526102
rect 21622 526046 21678 526102
rect 21250 525922 21306 525978
rect 21374 525922 21430 525978
rect 21498 525922 21554 525978
rect 21622 525922 21678 525978
rect 24970 598116 25026 598172
rect 25094 598116 25150 598172
rect 25218 598116 25274 598172
rect 25342 598116 25398 598172
rect 24970 597992 25026 598048
rect 25094 597992 25150 598048
rect 25218 597992 25274 598048
rect 25342 597992 25398 598048
rect 24970 597868 25026 597924
rect 25094 597868 25150 597924
rect 25218 597868 25274 597924
rect 25342 597868 25398 597924
rect 24970 597744 25026 597800
rect 25094 597744 25150 597800
rect 25218 597744 25274 597800
rect 25342 597744 25398 597800
rect 24970 586294 25026 586350
rect 25094 586294 25150 586350
rect 25218 586294 25274 586350
rect 25342 586294 25398 586350
rect 24970 586170 25026 586226
rect 25094 586170 25150 586226
rect 25218 586170 25274 586226
rect 25342 586170 25398 586226
rect 24970 586046 25026 586102
rect 25094 586046 25150 586102
rect 25218 586046 25274 586102
rect 25342 586046 25398 586102
rect 24970 585922 25026 585978
rect 25094 585922 25150 585978
rect 25218 585922 25274 585978
rect 25342 585922 25398 585978
rect 24970 568294 25026 568350
rect 25094 568294 25150 568350
rect 25218 568294 25274 568350
rect 25342 568294 25398 568350
rect 24970 568170 25026 568226
rect 25094 568170 25150 568226
rect 25218 568170 25274 568226
rect 25342 568170 25398 568226
rect 24970 568046 25026 568102
rect 25094 568046 25150 568102
rect 25218 568046 25274 568102
rect 25342 568046 25398 568102
rect 24970 567922 25026 567978
rect 25094 567922 25150 567978
rect 25218 567922 25274 567978
rect 25342 567922 25398 567978
rect 24970 550294 25026 550350
rect 25094 550294 25150 550350
rect 25218 550294 25274 550350
rect 25342 550294 25398 550350
rect 24970 550170 25026 550226
rect 25094 550170 25150 550226
rect 25218 550170 25274 550226
rect 25342 550170 25398 550226
rect 24970 550046 25026 550102
rect 25094 550046 25150 550102
rect 25218 550046 25274 550102
rect 25342 550046 25398 550102
rect 24970 549922 25026 549978
rect 25094 549922 25150 549978
rect 25218 549922 25274 549978
rect 25342 549922 25398 549978
rect 24970 532294 25026 532350
rect 25094 532294 25150 532350
rect 25218 532294 25274 532350
rect 25342 532294 25398 532350
rect 24970 532170 25026 532226
rect 25094 532170 25150 532226
rect 25218 532170 25274 532226
rect 25342 532170 25398 532226
rect 24970 532046 25026 532102
rect 25094 532046 25150 532102
rect 25218 532046 25274 532102
rect 25342 532046 25398 532102
rect 24970 531922 25026 531978
rect 25094 531922 25150 531978
rect 25218 531922 25274 531978
rect 25342 531922 25398 531978
rect 39250 597156 39306 597212
rect 39374 597156 39430 597212
rect 39498 597156 39554 597212
rect 39622 597156 39678 597212
rect 39250 597032 39306 597088
rect 39374 597032 39430 597088
rect 39498 597032 39554 597088
rect 39622 597032 39678 597088
rect 39250 596908 39306 596964
rect 39374 596908 39430 596964
rect 39498 596908 39554 596964
rect 39622 596908 39678 596964
rect 39250 596784 39306 596840
rect 39374 596784 39430 596840
rect 39498 596784 39554 596840
rect 39622 596784 39678 596840
rect 39250 580294 39306 580350
rect 39374 580294 39430 580350
rect 39498 580294 39554 580350
rect 39622 580294 39678 580350
rect 39250 580170 39306 580226
rect 39374 580170 39430 580226
rect 39498 580170 39554 580226
rect 39622 580170 39678 580226
rect 39250 580046 39306 580102
rect 39374 580046 39430 580102
rect 39498 580046 39554 580102
rect 39622 580046 39678 580102
rect 39250 579922 39306 579978
rect 39374 579922 39430 579978
rect 39498 579922 39554 579978
rect 39622 579922 39678 579978
rect 39250 562294 39306 562350
rect 39374 562294 39430 562350
rect 39498 562294 39554 562350
rect 39622 562294 39678 562350
rect 39250 562170 39306 562226
rect 39374 562170 39430 562226
rect 39498 562170 39554 562226
rect 39622 562170 39678 562226
rect 39250 562046 39306 562102
rect 39374 562046 39430 562102
rect 39498 562046 39554 562102
rect 39622 562046 39678 562102
rect 39250 561922 39306 561978
rect 39374 561922 39430 561978
rect 39498 561922 39554 561978
rect 39622 561922 39678 561978
rect 39250 544294 39306 544350
rect 39374 544294 39430 544350
rect 39498 544294 39554 544350
rect 39622 544294 39678 544350
rect 39250 544170 39306 544226
rect 39374 544170 39430 544226
rect 39498 544170 39554 544226
rect 39622 544170 39678 544226
rect 39250 544046 39306 544102
rect 39374 544046 39430 544102
rect 39498 544046 39554 544102
rect 39622 544046 39678 544102
rect 39250 543922 39306 543978
rect 39374 543922 39430 543978
rect 39498 543922 39554 543978
rect 39622 543922 39678 543978
rect 39250 526294 39306 526350
rect 39374 526294 39430 526350
rect 39498 526294 39554 526350
rect 39622 526294 39678 526350
rect 39250 526170 39306 526226
rect 39374 526170 39430 526226
rect 39498 526170 39554 526226
rect 39622 526170 39678 526226
rect 39250 526046 39306 526102
rect 39374 526046 39430 526102
rect 39498 526046 39554 526102
rect 39622 526046 39678 526102
rect 39250 525922 39306 525978
rect 39374 525922 39430 525978
rect 39498 525922 39554 525978
rect 39622 525922 39678 525978
rect 42970 598116 43026 598172
rect 43094 598116 43150 598172
rect 43218 598116 43274 598172
rect 43342 598116 43398 598172
rect 42970 597992 43026 598048
rect 43094 597992 43150 598048
rect 43218 597992 43274 598048
rect 43342 597992 43398 598048
rect 42970 597868 43026 597924
rect 43094 597868 43150 597924
rect 43218 597868 43274 597924
rect 43342 597868 43398 597924
rect 42970 597744 43026 597800
rect 43094 597744 43150 597800
rect 43218 597744 43274 597800
rect 43342 597744 43398 597800
rect 42970 586294 43026 586350
rect 43094 586294 43150 586350
rect 43218 586294 43274 586350
rect 43342 586294 43398 586350
rect 42970 586170 43026 586226
rect 43094 586170 43150 586226
rect 43218 586170 43274 586226
rect 43342 586170 43398 586226
rect 42970 586046 43026 586102
rect 43094 586046 43150 586102
rect 43218 586046 43274 586102
rect 43342 586046 43398 586102
rect 42970 585922 43026 585978
rect 43094 585922 43150 585978
rect 43218 585922 43274 585978
rect 43342 585922 43398 585978
rect 42970 568294 43026 568350
rect 43094 568294 43150 568350
rect 43218 568294 43274 568350
rect 43342 568294 43398 568350
rect 42970 568170 43026 568226
rect 43094 568170 43150 568226
rect 43218 568170 43274 568226
rect 43342 568170 43398 568226
rect 42970 568046 43026 568102
rect 43094 568046 43150 568102
rect 43218 568046 43274 568102
rect 43342 568046 43398 568102
rect 42970 567922 43026 567978
rect 43094 567922 43150 567978
rect 43218 567922 43274 567978
rect 43342 567922 43398 567978
rect 42970 550294 43026 550350
rect 43094 550294 43150 550350
rect 43218 550294 43274 550350
rect 43342 550294 43398 550350
rect 42970 550170 43026 550226
rect 43094 550170 43150 550226
rect 43218 550170 43274 550226
rect 43342 550170 43398 550226
rect 42970 550046 43026 550102
rect 43094 550046 43150 550102
rect 43218 550046 43274 550102
rect 43342 550046 43398 550102
rect 42970 549922 43026 549978
rect 43094 549922 43150 549978
rect 43218 549922 43274 549978
rect 43342 549922 43398 549978
rect 42970 532294 43026 532350
rect 43094 532294 43150 532350
rect 43218 532294 43274 532350
rect 43342 532294 43398 532350
rect 42970 532170 43026 532226
rect 43094 532170 43150 532226
rect 43218 532170 43274 532226
rect 43342 532170 43398 532226
rect 42970 532046 43026 532102
rect 43094 532046 43150 532102
rect 43218 532046 43274 532102
rect 43342 532046 43398 532102
rect 42970 531922 43026 531978
rect 43094 531922 43150 531978
rect 43218 531922 43274 531978
rect 43342 531922 43398 531978
rect 57250 597156 57306 597212
rect 57374 597156 57430 597212
rect 57498 597156 57554 597212
rect 57622 597156 57678 597212
rect 57250 597032 57306 597088
rect 57374 597032 57430 597088
rect 57498 597032 57554 597088
rect 57622 597032 57678 597088
rect 57250 596908 57306 596964
rect 57374 596908 57430 596964
rect 57498 596908 57554 596964
rect 57622 596908 57678 596964
rect 57250 596784 57306 596840
rect 57374 596784 57430 596840
rect 57498 596784 57554 596840
rect 57622 596784 57678 596840
rect 57250 580294 57306 580350
rect 57374 580294 57430 580350
rect 57498 580294 57554 580350
rect 57622 580294 57678 580350
rect 57250 580170 57306 580226
rect 57374 580170 57430 580226
rect 57498 580170 57554 580226
rect 57622 580170 57678 580226
rect 57250 580046 57306 580102
rect 57374 580046 57430 580102
rect 57498 580046 57554 580102
rect 57622 580046 57678 580102
rect 57250 579922 57306 579978
rect 57374 579922 57430 579978
rect 57498 579922 57554 579978
rect 57622 579922 57678 579978
rect 57250 562294 57306 562350
rect 57374 562294 57430 562350
rect 57498 562294 57554 562350
rect 57622 562294 57678 562350
rect 57250 562170 57306 562226
rect 57374 562170 57430 562226
rect 57498 562170 57554 562226
rect 57622 562170 57678 562226
rect 57250 562046 57306 562102
rect 57374 562046 57430 562102
rect 57498 562046 57554 562102
rect 57622 562046 57678 562102
rect 57250 561922 57306 561978
rect 57374 561922 57430 561978
rect 57498 561922 57554 561978
rect 57622 561922 57678 561978
rect 57250 544294 57306 544350
rect 57374 544294 57430 544350
rect 57498 544294 57554 544350
rect 57622 544294 57678 544350
rect 57250 544170 57306 544226
rect 57374 544170 57430 544226
rect 57498 544170 57554 544226
rect 57622 544170 57678 544226
rect 57250 544046 57306 544102
rect 57374 544046 57430 544102
rect 57498 544046 57554 544102
rect 57622 544046 57678 544102
rect 57250 543922 57306 543978
rect 57374 543922 57430 543978
rect 57498 543922 57554 543978
rect 57622 543922 57678 543978
rect 57250 526294 57306 526350
rect 57374 526294 57430 526350
rect 57498 526294 57554 526350
rect 57622 526294 57678 526350
rect 57250 526170 57306 526226
rect 57374 526170 57430 526226
rect 57498 526170 57554 526226
rect 57622 526170 57678 526226
rect 57250 526046 57306 526102
rect 57374 526046 57430 526102
rect 57498 526046 57554 526102
rect 57622 526046 57678 526102
rect 57250 525922 57306 525978
rect 57374 525922 57430 525978
rect 57498 525922 57554 525978
rect 57622 525922 57678 525978
rect 60970 598116 61026 598172
rect 61094 598116 61150 598172
rect 61218 598116 61274 598172
rect 61342 598116 61398 598172
rect 60970 597992 61026 598048
rect 61094 597992 61150 598048
rect 61218 597992 61274 598048
rect 61342 597992 61398 598048
rect 60970 597868 61026 597924
rect 61094 597868 61150 597924
rect 61218 597868 61274 597924
rect 61342 597868 61398 597924
rect 60970 597744 61026 597800
rect 61094 597744 61150 597800
rect 61218 597744 61274 597800
rect 61342 597744 61398 597800
rect 60970 586294 61026 586350
rect 61094 586294 61150 586350
rect 61218 586294 61274 586350
rect 61342 586294 61398 586350
rect 60970 586170 61026 586226
rect 61094 586170 61150 586226
rect 61218 586170 61274 586226
rect 61342 586170 61398 586226
rect 60970 586046 61026 586102
rect 61094 586046 61150 586102
rect 61218 586046 61274 586102
rect 61342 586046 61398 586102
rect 60970 585922 61026 585978
rect 61094 585922 61150 585978
rect 61218 585922 61274 585978
rect 61342 585922 61398 585978
rect 60970 568294 61026 568350
rect 61094 568294 61150 568350
rect 61218 568294 61274 568350
rect 61342 568294 61398 568350
rect 60970 568170 61026 568226
rect 61094 568170 61150 568226
rect 61218 568170 61274 568226
rect 61342 568170 61398 568226
rect 60970 568046 61026 568102
rect 61094 568046 61150 568102
rect 61218 568046 61274 568102
rect 61342 568046 61398 568102
rect 60970 567922 61026 567978
rect 61094 567922 61150 567978
rect 61218 567922 61274 567978
rect 61342 567922 61398 567978
rect 60970 550294 61026 550350
rect 61094 550294 61150 550350
rect 61218 550294 61274 550350
rect 61342 550294 61398 550350
rect 60970 550170 61026 550226
rect 61094 550170 61150 550226
rect 61218 550170 61274 550226
rect 61342 550170 61398 550226
rect 60970 550046 61026 550102
rect 61094 550046 61150 550102
rect 61218 550046 61274 550102
rect 61342 550046 61398 550102
rect 60970 549922 61026 549978
rect 61094 549922 61150 549978
rect 61218 549922 61274 549978
rect 61342 549922 61398 549978
rect 60970 532294 61026 532350
rect 61094 532294 61150 532350
rect 61218 532294 61274 532350
rect 61342 532294 61398 532350
rect 60970 532170 61026 532226
rect 61094 532170 61150 532226
rect 61218 532170 61274 532226
rect 61342 532170 61398 532226
rect 60970 532046 61026 532102
rect 61094 532046 61150 532102
rect 61218 532046 61274 532102
rect 61342 532046 61398 532102
rect 60970 531922 61026 531978
rect 61094 531922 61150 531978
rect 61218 531922 61274 531978
rect 61342 531922 61398 531978
rect 75250 597156 75306 597212
rect 75374 597156 75430 597212
rect 75498 597156 75554 597212
rect 75622 597156 75678 597212
rect 75250 597032 75306 597088
rect 75374 597032 75430 597088
rect 75498 597032 75554 597088
rect 75622 597032 75678 597088
rect 75250 596908 75306 596964
rect 75374 596908 75430 596964
rect 75498 596908 75554 596964
rect 75622 596908 75678 596964
rect 75250 596784 75306 596840
rect 75374 596784 75430 596840
rect 75498 596784 75554 596840
rect 75622 596784 75678 596840
rect 75250 580294 75306 580350
rect 75374 580294 75430 580350
rect 75498 580294 75554 580350
rect 75622 580294 75678 580350
rect 75250 580170 75306 580226
rect 75374 580170 75430 580226
rect 75498 580170 75554 580226
rect 75622 580170 75678 580226
rect 75250 580046 75306 580102
rect 75374 580046 75430 580102
rect 75498 580046 75554 580102
rect 75622 580046 75678 580102
rect 75250 579922 75306 579978
rect 75374 579922 75430 579978
rect 75498 579922 75554 579978
rect 75622 579922 75678 579978
rect 75250 562294 75306 562350
rect 75374 562294 75430 562350
rect 75498 562294 75554 562350
rect 75622 562294 75678 562350
rect 75250 562170 75306 562226
rect 75374 562170 75430 562226
rect 75498 562170 75554 562226
rect 75622 562170 75678 562226
rect 75250 562046 75306 562102
rect 75374 562046 75430 562102
rect 75498 562046 75554 562102
rect 75622 562046 75678 562102
rect 75250 561922 75306 561978
rect 75374 561922 75430 561978
rect 75498 561922 75554 561978
rect 75622 561922 75678 561978
rect 75250 544294 75306 544350
rect 75374 544294 75430 544350
rect 75498 544294 75554 544350
rect 75622 544294 75678 544350
rect 75250 544170 75306 544226
rect 75374 544170 75430 544226
rect 75498 544170 75554 544226
rect 75622 544170 75678 544226
rect 75250 544046 75306 544102
rect 75374 544046 75430 544102
rect 75498 544046 75554 544102
rect 75622 544046 75678 544102
rect 75250 543922 75306 543978
rect 75374 543922 75430 543978
rect 75498 543922 75554 543978
rect 75622 543922 75678 543978
rect 75250 526294 75306 526350
rect 75374 526294 75430 526350
rect 75498 526294 75554 526350
rect 75622 526294 75678 526350
rect 75250 526170 75306 526226
rect 75374 526170 75430 526226
rect 75498 526170 75554 526226
rect 75622 526170 75678 526226
rect 75250 526046 75306 526102
rect 75374 526046 75430 526102
rect 75498 526046 75554 526102
rect 75622 526046 75678 526102
rect 75250 525922 75306 525978
rect 75374 525922 75430 525978
rect 75498 525922 75554 525978
rect 75622 525922 75678 525978
rect 78970 598116 79026 598172
rect 79094 598116 79150 598172
rect 79218 598116 79274 598172
rect 79342 598116 79398 598172
rect 78970 597992 79026 598048
rect 79094 597992 79150 598048
rect 79218 597992 79274 598048
rect 79342 597992 79398 598048
rect 78970 597868 79026 597924
rect 79094 597868 79150 597924
rect 79218 597868 79274 597924
rect 79342 597868 79398 597924
rect 78970 597744 79026 597800
rect 79094 597744 79150 597800
rect 79218 597744 79274 597800
rect 79342 597744 79398 597800
rect 78970 586294 79026 586350
rect 79094 586294 79150 586350
rect 79218 586294 79274 586350
rect 79342 586294 79398 586350
rect 78970 586170 79026 586226
rect 79094 586170 79150 586226
rect 79218 586170 79274 586226
rect 79342 586170 79398 586226
rect 78970 586046 79026 586102
rect 79094 586046 79150 586102
rect 79218 586046 79274 586102
rect 79342 586046 79398 586102
rect 78970 585922 79026 585978
rect 79094 585922 79150 585978
rect 79218 585922 79274 585978
rect 79342 585922 79398 585978
rect 78970 568294 79026 568350
rect 79094 568294 79150 568350
rect 79218 568294 79274 568350
rect 79342 568294 79398 568350
rect 78970 568170 79026 568226
rect 79094 568170 79150 568226
rect 79218 568170 79274 568226
rect 79342 568170 79398 568226
rect 78970 568046 79026 568102
rect 79094 568046 79150 568102
rect 79218 568046 79274 568102
rect 79342 568046 79398 568102
rect 78970 567922 79026 567978
rect 79094 567922 79150 567978
rect 79218 567922 79274 567978
rect 79342 567922 79398 567978
rect 78970 550294 79026 550350
rect 79094 550294 79150 550350
rect 79218 550294 79274 550350
rect 79342 550294 79398 550350
rect 78970 550170 79026 550226
rect 79094 550170 79150 550226
rect 79218 550170 79274 550226
rect 79342 550170 79398 550226
rect 78970 550046 79026 550102
rect 79094 550046 79150 550102
rect 79218 550046 79274 550102
rect 79342 550046 79398 550102
rect 78970 549922 79026 549978
rect 79094 549922 79150 549978
rect 79218 549922 79274 549978
rect 79342 549922 79398 549978
rect 78970 532294 79026 532350
rect 79094 532294 79150 532350
rect 79218 532294 79274 532350
rect 79342 532294 79398 532350
rect 78970 532170 79026 532226
rect 79094 532170 79150 532226
rect 79218 532170 79274 532226
rect 79342 532170 79398 532226
rect 78970 532046 79026 532102
rect 79094 532046 79150 532102
rect 79218 532046 79274 532102
rect 79342 532046 79398 532102
rect 78970 531922 79026 531978
rect 79094 531922 79150 531978
rect 79218 531922 79274 531978
rect 79342 531922 79398 531978
rect 93250 597156 93306 597212
rect 93374 597156 93430 597212
rect 93498 597156 93554 597212
rect 93622 597156 93678 597212
rect 93250 597032 93306 597088
rect 93374 597032 93430 597088
rect 93498 597032 93554 597088
rect 93622 597032 93678 597088
rect 93250 596908 93306 596964
rect 93374 596908 93430 596964
rect 93498 596908 93554 596964
rect 93622 596908 93678 596964
rect 93250 596784 93306 596840
rect 93374 596784 93430 596840
rect 93498 596784 93554 596840
rect 93622 596784 93678 596840
rect 93250 580294 93306 580350
rect 93374 580294 93430 580350
rect 93498 580294 93554 580350
rect 93622 580294 93678 580350
rect 93250 580170 93306 580226
rect 93374 580170 93430 580226
rect 93498 580170 93554 580226
rect 93622 580170 93678 580226
rect 93250 580046 93306 580102
rect 93374 580046 93430 580102
rect 93498 580046 93554 580102
rect 93622 580046 93678 580102
rect 93250 579922 93306 579978
rect 93374 579922 93430 579978
rect 93498 579922 93554 579978
rect 93622 579922 93678 579978
rect 93250 562294 93306 562350
rect 93374 562294 93430 562350
rect 93498 562294 93554 562350
rect 93622 562294 93678 562350
rect 93250 562170 93306 562226
rect 93374 562170 93430 562226
rect 93498 562170 93554 562226
rect 93622 562170 93678 562226
rect 93250 562046 93306 562102
rect 93374 562046 93430 562102
rect 93498 562046 93554 562102
rect 93622 562046 93678 562102
rect 93250 561922 93306 561978
rect 93374 561922 93430 561978
rect 93498 561922 93554 561978
rect 93622 561922 93678 561978
rect 93250 544294 93306 544350
rect 93374 544294 93430 544350
rect 93498 544294 93554 544350
rect 93622 544294 93678 544350
rect 93250 544170 93306 544226
rect 93374 544170 93430 544226
rect 93498 544170 93554 544226
rect 93622 544170 93678 544226
rect 93250 544046 93306 544102
rect 93374 544046 93430 544102
rect 93498 544046 93554 544102
rect 93622 544046 93678 544102
rect 93250 543922 93306 543978
rect 93374 543922 93430 543978
rect 93498 543922 93554 543978
rect 93622 543922 93678 543978
rect 93250 526294 93306 526350
rect 93374 526294 93430 526350
rect 93498 526294 93554 526350
rect 93622 526294 93678 526350
rect 93250 526170 93306 526226
rect 93374 526170 93430 526226
rect 93498 526170 93554 526226
rect 93622 526170 93678 526226
rect 93250 526046 93306 526102
rect 93374 526046 93430 526102
rect 93498 526046 93554 526102
rect 93622 526046 93678 526102
rect 93250 525922 93306 525978
rect 93374 525922 93430 525978
rect 93498 525922 93554 525978
rect 93622 525922 93678 525978
rect 96970 598116 97026 598172
rect 97094 598116 97150 598172
rect 97218 598116 97274 598172
rect 97342 598116 97398 598172
rect 96970 597992 97026 598048
rect 97094 597992 97150 598048
rect 97218 597992 97274 598048
rect 97342 597992 97398 598048
rect 96970 597868 97026 597924
rect 97094 597868 97150 597924
rect 97218 597868 97274 597924
rect 97342 597868 97398 597924
rect 96970 597744 97026 597800
rect 97094 597744 97150 597800
rect 97218 597744 97274 597800
rect 97342 597744 97398 597800
rect 96970 586294 97026 586350
rect 97094 586294 97150 586350
rect 97218 586294 97274 586350
rect 97342 586294 97398 586350
rect 96970 586170 97026 586226
rect 97094 586170 97150 586226
rect 97218 586170 97274 586226
rect 97342 586170 97398 586226
rect 96970 586046 97026 586102
rect 97094 586046 97150 586102
rect 97218 586046 97274 586102
rect 97342 586046 97398 586102
rect 96970 585922 97026 585978
rect 97094 585922 97150 585978
rect 97218 585922 97274 585978
rect 97342 585922 97398 585978
rect 96970 568294 97026 568350
rect 97094 568294 97150 568350
rect 97218 568294 97274 568350
rect 97342 568294 97398 568350
rect 96970 568170 97026 568226
rect 97094 568170 97150 568226
rect 97218 568170 97274 568226
rect 97342 568170 97398 568226
rect 96970 568046 97026 568102
rect 97094 568046 97150 568102
rect 97218 568046 97274 568102
rect 97342 568046 97398 568102
rect 96970 567922 97026 567978
rect 97094 567922 97150 567978
rect 97218 567922 97274 567978
rect 97342 567922 97398 567978
rect 96970 550294 97026 550350
rect 97094 550294 97150 550350
rect 97218 550294 97274 550350
rect 97342 550294 97398 550350
rect 96970 550170 97026 550226
rect 97094 550170 97150 550226
rect 97218 550170 97274 550226
rect 97342 550170 97398 550226
rect 96970 550046 97026 550102
rect 97094 550046 97150 550102
rect 97218 550046 97274 550102
rect 97342 550046 97398 550102
rect 96970 549922 97026 549978
rect 97094 549922 97150 549978
rect 97218 549922 97274 549978
rect 97342 549922 97398 549978
rect 96970 532294 97026 532350
rect 97094 532294 97150 532350
rect 97218 532294 97274 532350
rect 97342 532294 97398 532350
rect 96970 532170 97026 532226
rect 97094 532170 97150 532226
rect 97218 532170 97274 532226
rect 97342 532170 97398 532226
rect 96970 532046 97026 532102
rect 97094 532046 97150 532102
rect 97218 532046 97274 532102
rect 97342 532046 97398 532102
rect 96970 531922 97026 531978
rect 97094 531922 97150 531978
rect 97218 531922 97274 531978
rect 97342 531922 97398 531978
rect 111250 597156 111306 597212
rect 111374 597156 111430 597212
rect 111498 597156 111554 597212
rect 111622 597156 111678 597212
rect 111250 597032 111306 597088
rect 111374 597032 111430 597088
rect 111498 597032 111554 597088
rect 111622 597032 111678 597088
rect 111250 596908 111306 596964
rect 111374 596908 111430 596964
rect 111498 596908 111554 596964
rect 111622 596908 111678 596964
rect 111250 596784 111306 596840
rect 111374 596784 111430 596840
rect 111498 596784 111554 596840
rect 111622 596784 111678 596840
rect 111250 580294 111306 580350
rect 111374 580294 111430 580350
rect 111498 580294 111554 580350
rect 111622 580294 111678 580350
rect 111250 580170 111306 580226
rect 111374 580170 111430 580226
rect 111498 580170 111554 580226
rect 111622 580170 111678 580226
rect 111250 580046 111306 580102
rect 111374 580046 111430 580102
rect 111498 580046 111554 580102
rect 111622 580046 111678 580102
rect 111250 579922 111306 579978
rect 111374 579922 111430 579978
rect 111498 579922 111554 579978
rect 111622 579922 111678 579978
rect 111250 562294 111306 562350
rect 111374 562294 111430 562350
rect 111498 562294 111554 562350
rect 111622 562294 111678 562350
rect 111250 562170 111306 562226
rect 111374 562170 111430 562226
rect 111498 562170 111554 562226
rect 111622 562170 111678 562226
rect 111250 562046 111306 562102
rect 111374 562046 111430 562102
rect 111498 562046 111554 562102
rect 111622 562046 111678 562102
rect 111250 561922 111306 561978
rect 111374 561922 111430 561978
rect 111498 561922 111554 561978
rect 111622 561922 111678 561978
rect 111250 544294 111306 544350
rect 111374 544294 111430 544350
rect 111498 544294 111554 544350
rect 111622 544294 111678 544350
rect 111250 544170 111306 544226
rect 111374 544170 111430 544226
rect 111498 544170 111554 544226
rect 111622 544170 111678 544226
rect 111250 544046 111306 544102
rect 111374 544046 111430 544102
rect 111498 544046 111554 544102
rect 111622 544046 111678 544102
rect 111250 543922 111306 543978
rect 111374 543922 111430 543978
rect 111498 543922 111554 543978
rect 111622 543922 111678 543978
rect 111250 526294 111306 526350
rect 111374 526294 111430 526350
rect 111498 526294 111554 526350
rect 111622 526294 111678 526350
rect 111250 526170 111306 526226
rect 111374 526170 111430 526226
rect 111498 526170 111554 526226
rect 111622 526170 111678 526226
rect 111250 526046 111306 526102
rect 111374 526046 111430 526102
rect 111498 526046 111554 526102
rect 111622 526046 111678 526102
rect 111250 525922 111306 525978
rect 111374 525922 111430 525978
rect 111498 525922 111554 525978
rect 111622 525922 111678 525978
rect 114970 598116 115026 598172
rect 115094 598116 115150 598172
rect 115218 598116 115274 598172
rect 115342 598116 115398 598172
rect 114970 597992 115026 598048
rect 115094 597992 115150 598048
rect 115218 597992 115274 598048
rect 115342 597992 115398 598048
rect 114970 597868 115026 597924
rect 115094 597868 115150 597924
rect 115218 597868 115274 597924
rect 115342 597868 115398 597924
rect 114970 597744 115026 597800
rect 115094 597744 115150 597800
rect 115218 597744 115274 597800
rect 115342 597744 115398 597800
rect 114970 586294 115026 586350
rect 115094 586294 115150 586350
rect 115218 586294 115274 586350
rect 115342 586294 115398 586350
rect 114970 586170 115026 586226
rect 115094 586170 115150 586226
rect 115218 586170 115274 586226
rect 115342 586170 115398 586226
rect 114970 586046 115026 586102
rect 115094 586046 115150 586102
rect 115218 586046 115274 586102
rect 115342 586046 115398 586102
rect 114970 585922 115026 585978
rect 115094 585922 115150 585978
rect 115218 585922 115274 585978
rect 115342 585922 115398 585978
rect 114970 568294 115026 568350
rect 115094 568294 115150 568350
rect 115218 568294 115274 568350
rect 115342 568294 115398 568350
rect 114970 568170 115026 568226
rect 115094 568170 115150 568226
rect 115218 568170 115274 568226
rect 115342 568170 115398 568226
rect 114970 568046 115026 568102
rect 115094 568046 115150 568102
rect 115218 568046 115274 568102
rect 115342 568046 115398 568102
rect 114970 567922 115026 567978
rect 115094 567922 115150 567978
rect 115218 567922 115274 567978
rect 115342 567922 115398 567978
rect 114970 550294 115026 550350
rect 115094 550294 115150 550350
rect 115218 550294 115274 550350
rect 115342 550294 115398 550350
rect 114970 550170 115026 550226
rect 115094 550170 115150 550226
rect 115218 550170 115274 550226
rect 115342 550170 115398 550226
rect 114970 550046 115026 550102
rect 115094 550046 115150 550102
rect 115218 550046 115274 550102
rect 115342 550046 115398 550102
rect 114970 549922 115026 549978
rect 115094 549922 115150 549978
rect 115218 549922 115274 549978
rect 115342 549922 115398 549978
rect 114970 532294 115026 532350
rect 115094 532294 115150 532350
rect 115218 532294 115274 532350
rect 115342 532294 115398 532350
rect 114970 532170 115026 532226
rect 115094 532170 115150 532226
rect 115218 532170 115274 532226
rect 115342 532170 115398 532226
rect 114970 532046 115026 532102
rect 115094 532046 115150 532102
rect 115218 532046 115274 532102
rect 115342 532046 115398 532102
rect 114970 531922 115026 531978
rect 115094 531922 115150 531978
rect 115218 531922 115274 531978
rect 115342 531922 115398 531978
rect 129250 597156 129306 597212
rect 129374 597156 129430 597212
rect 129498 597156 129554 597212
rect 129622 597156 129678 597212
rect 129250 597032 129306 597088
rect 129374 597032 129430 597088
rect 129498 597032 129554 597088
rect 129622 597032 129678 597088
rect 129250 596908 129306 596964
rect 129374 596908 129430 596964
rect 129498 596908 129554 596964
rect 129622 596908 129678 596964
rect 129250 596784 129306 596840
rect 129374 596784 129430 596840
rect 129498 596784 129554 596840
rect 129622 596784 129678 596840
rect 129250 580294 129306 580350
rect 129374 580294 129430 580350
rect 129498 580294 129554 580350
rect 129622 580294 129678 580350
rect 129250 580170 129306 580226
rect 129374 580170 129430 580226
rect 129498 580170 129554 580226
rect 129622 580170 129678 580226
rect 129250 580046 129306 580102
rect 129374 580046 129430 580102
rect 129498 580046 129554 580102
rect 129622 580046 129678 580102
rect 129250 579922 129306 579978
rect 129374 579922 129430 579978
rect 129498 579922 129554 579978
rect 129622 579922 129678 579978
rect 129250 562294 129306 562350
rect 129374 562294 129430 562350
rect 129498 562294 129554 562350
rect 129622 562294 129678 562350
rect 129250 562170 129306 562226
rect 129374 562170 129430 562226
rect 129498 562170 129554 562226
rect 129622 562170 129678 562226
rect 129250 562046 129306 562102
rect 129374 562046 129430 562102
rect 129498 562046 129554 562102
rect 129622 562046 129678 562102
rect 129250 561922 129306 561978
rect 129374 561922 129430 561978
rect 129498 561922 129554 561978
rect 129622 561922 129678 561978
rect 129250 544294 129306 544350
rect 129374 544294 129430 544350
rect 129498 544294 129554 544350
rect 129622 544294 129678 544350
rect 129250 544170 129306 544226
rect 129374 544170 129430 544226
rect 129498 544170 129554 544226
rect 129622 544170 129678 544226
rect 129250 544046 129306 544102
rect 129374 544046 129430 544102
rect 129498 544046 129554 544102
rect 129622 544046 129678 544102
rect 129250 543922 129306 543978
rect 129374 543922 129430 543978
rect 129498 543922 129554 543978
rect 129622 543922 129678 543978
rect 129250 526294 129306 526350
rect 129374 526294 129430 526350
rect 129498 526294 129554 526350
rect 129622 526294 129678 526350
rect 129250 526170 129306 526226
rect 129374 526170 129430 526226
rect 129498 526170 129554 526226
rect 129622 526170 129678 526226
rect 129250 526046 129306 526102
rect 129374 526046 129430 526102
rect 129498 526046 129554 526102
rect 129622 526046 129678 526102
rect 129250 525922 129306 525978
rect 129374 525922 129430 525978
rect 129498 525922 129554 525978
rect 129622 525922 129678 525978
rect 132970 598116 133026 598172
rect 133094 598116 133150 598172
rect 133218 598116 133274 598172
rect 133342 598116 133398 598172
rect 132970 597992 133026 598048
rect 133094 597992 133150 598048
rect 133218 597992 133274 598048
rect 133342 597992 133398 598048
rect 132970 597868 133026 597924
rect 133094 597868 133150 597924
rect 133218 597868 133274 597924
rect 133342 597868 133398 597924
rect 132970 597744 133026 597800
rect 133094 597744 133150 597800
rect 133218 597744 133274 597800
rect 133342 597744 133398 597800
rect 132970 586294 133026 586350
rect 133094 586294 133150 586350
rect 133218 586294 133274 586350
rect 133342 586294 133398 586350
rect 132970 586170 133026 586226
rect 133094 586170 133150 586226
rect 133218 586170 133274 586226
rect 133342 586170 133398 586226
rect 132970 586046 133026 586102
rect 133094 586046 133150 586102
rect 133218 586046 133274 586102
rect 133342 586046 133398 586102
rect 132970 585922 133026 585978
rect 133094 585922 133150 585978
rect 133218 585922 133274 585978
rect 133342 585922 133398 585978
rect 132970 568294 133026 568350
rect 133094 568294 133150 568350
rect 133218 568294 133274 568350
rect 133342 568294 133398 568350
rect 132970 568170 133026 568226
rect 133094 568170 133150 568226
rect 133218 568170 133274 568226
rect 133342 568170 133398 568226
rect 132970 568046 133026 568102
rect 133094 568046 133150 568102
rect 133218 568046 133274 568102
rect 133342 568046 133398 568102
rect 132970 567922 133026 567978
rect 133094 567922 133150 567978
rect 133218 567922 133274 567978
rect 133342 567922 133398 567978
rect 132970 550294 133026 550350
rect 133094 550294 133150 550350
rect 133218 550294 133274 550350
rect 133342 550294 133398 550350
rect 132970 550170 133026 550226
rect 133094 550170 133150 550226
rect 133218 550170 133274 550226
rect 133342 550170 133398 550226
rect 132970 550046 133026 550102
rect 133094 550046 133150 550102
rect 133218 550046 133274 550102
rect 133342 550046 133398 550102
rect 132970 549922 133026 549978
rect 133094 549922 133150 549978
rect 133218 549922 133274 549978
rect 133342 549922 133398 549978
rect 132970 532294 133026 532350
rect 133094 532294 133150 532350
rect 133218 532294 133274 532350
rect 133342 532294 133398 532350
rect 132970 532170 133026 532226
rect 133094 532170 133150 532226
rect 133218 532170 133274 532226
rect 133342 532170 133398 532226
rect 132970 532046 133026 532102
rect 133094 532046 133150 532102
rect 133218 532046 133274 532102
rect 133342 532046 133398 532102
rect 132970 531922 133026 531978
rect 133094 531922 133150 531978
rect 133218 531922 133274 531978
rect 133342 531922 133398 531978
rect 147250 597156 147306 597212
rect 147374 597156 147430 597212
rect 147498 597156 147554 597212
rect 147622 597156 147678 597212
rect 147250 597032 147306 597088
rect 147374 597032 147430 597088
rect 147498 597032 147554 597088
rect 147622 597032 147678 597088
rect 147250 596908 147306 596964
rect 147374 596908 147430 596964
rect 147498 596908 147554 596964
rect 147622 596908 147678 596964
rect 147250 596784 147306 596840
rect 147374 596784 147430 596840
rect 147498 596784 147554 596840
rect 147622 596784 147678 596840
rect 147250 580294 147306 580350
rect 147374 580294 147430 580350
rect 147498 580294 147554 580350
rect 147622 580294 147678 580350
rect 147250 580170 147306 580226
rect 147374 580170 147430 580226
rect 147498 580170 147554 580226
rect 147622 580170 147678 580226
rect 147250 580046 147306 580102
rect 147374 580046 147430 580102
rect 147498 580046 147554 580102
rect 147622 580046 147678 580102
rect 147250 579922 147306 579978
rect 147374 579922 147430 579978
rect 147498 579922 147554 579978
rect 147622 579922 147678 579978
rect 147250 562294 147306 562350
rect 147374 562294 147430 562350
rect 147498 562294 147554 562350
rect 147622 562294 147678 562350
rect 147250 562170 147306 562226
rect 147374 562170 147430 562226
rect 147498 562170 147554 562226
rect 147622 562170 147678 562226
rect 147250 562046 147306 562102
rect 147374 562046 147430 562102
rect 147498 562046 147554 562102
rect 147622 562046 147678 562102
rect 147250 561922 147306 561978
rect 147374 561922 147430 561978
rect 147498 561922 147554 561978
rect 147622 561922 147678 561978
rect 147250 544294 147306 544350
rect 147374 544294 147430 544350
rect 147498 544294 147554 544350
rect 147622 544294 147678 544350
rect 147250 544170 147306 544226
rect 147374 544170 147430 544226
rect 147498 544170 147554 544226
rect 147622 544170 147678 544226
rect 147250 544046 147306 544102
rect 147374 544046 147430 544102
rect 147498 544046 147554 544102
rect 147622 544046 147678 544102
rect 147250 543922 147306 543978
rect 147374 543922 147430 543978
rect 147498 543922 147554 543978
rect 147622 543922 147678 543978
rect 147250 526294 147306 526350
rect 147374 526294 147430 526350
rect 147498 526294 147554 526350
rect 147622 526294 147678 526350
rect 147250 526170 147306 526226
rect 147374 526170 147430 526226
rect 147498 526170 147554 526226
rect 147622 526170 147678 526226
rect 147250 526046 147306 526102
rect 147374 526046 147430 526102
rect 147498 526046 147554 526102
rect 147622 526046 147678 526102
rect 147250 525922 147306 525978
rect 147374 525922 147430 525978
rect 147498 525922 147554 525978
rect 147622 525922 147678 525978
rect 150970 598116 151026 598172
rect 151094 598116 151150 598172
rect 151218 598116 151274 598172
rect 151342 598116 151398 598172
rect 150970 597992 151026 598048
rect 151094 597992 151150 598048
rect 151218 597992 151274 598048
rect 151342 597992 151398 598048
rect 150970 597868 151026 597924
rect 151094 597868 151150 597924
rect 151218 597868 151274 597924
rect 151342 597868 151398 597924
rect 150970 597744 151026 597800
rect 151094 597744 151150 597800
rect 151218 597744 151274 597800
rect 151342 597744 151398 597800
rect 150970 586294 151026 586350
rect 151094 586294 151150 586350
rect 151218 586294 151274 586350
rect 151342 586294 151398 586350
rect 150970 586170 151026 586226
rect 151094 586170 151150 586226
rect 151218 586170 151274 586226
rect 151342 586170 151398 586226
rect 150970 586046 151026 586102
rect 151094 586046 151150 586102
rect 151218 586046 151274 586102
rect 151342 586046 151398 586102
rect 150970 585922 151026 585978
rect 151094 585922 151150 585978
rect 151218 585922 151274 585978
rect 151342 585922 151398 585978
rect 150970 568294 151026 568350
rect 151094 568294 151150 568350
rect 151218 568294 151274 568350
rect 151342 568294 151398 568350
rect 150970 568170 151026 568226
rect 151094 568170 151150 568226
rect 151218 568170 151274 568226
rect 151342 568170 151398 568226
rect 150970 568046 151026 568102
rect 151094 568046 151150 568102
rect 151218 568046 151274 568102
rect 151342 568046 151398 568102
rect 150970 567922 151026 567978
rect 151094 567922 151150 567978
rect 151218 567922 151274 567978
rect 151342 567922 151398 567978
rect 150970 550294 151026 550350
rect 151094 550294 151150 550350
rect 151218 550294 151274 550350
rect 151342 550294 151398 550350
rect 150970 550170 151026 550226
rect 151094 550170 151150 550226
rect 151218 550170 151274 550226
rect 151342 550170 151398 550226
rect 150970 550046 151026 550102
rect 151094 550046 151150 550102
rect 151218 550046 151274 550102
rect 151342 550046 151398 550102
rect 150970 549922 151026 549978
rect 151094 549922 151150 549978
rect 151218 549922 151274 549978
rect 151342 549922 151398 549978
rect 150970 532294 151026 532350
rect 151094 532294 151150 532350
rect 151218 532294 151274 532350
rect 151342 532294 151398 532350
rect 150970 532170 151026 532226
rect 151094 532170 151150 532226
rect 151218 532170 151274 532226
rect 151342 532170 151398 532226
rect 150970 532046 151026 532102
rect 151094 532046 151150 532102
rect 151218 532046 151274 532102
rect 151342 532046 151398 532102
rect 150970 531922 151026 531978
rect 151094 531922 151150 531978
rect 151218 531922 151274 531978
rect 151342 531922 151398 531978
rect 165250 597156 165306 597212
rect 165374 597156 165430 597212
rect 165498 597156 165554 597212
rect 165622 597156 165678 597212
rect 165250 597032 165306 597088
rect 165374 597032 165430 597088
rect 165498 597032 165554 597088
rect 165622 597032 165678 597088
rect 165250 596908 165306 596964
rect 165374 596908 165430 596964
rect 165498 596908 165554 596964
rect 165622 596908 165678 596964
rect 165250 596784 165306 596840
rect 165374 596784 165430 596840
rect 165498 596784 165554 596840
rect 165622 596784 165678 596840
rect 165250 580294 165306 580350
rect 165374 580294 165430 580350
rect 165498 580294 165554 580350
rect 165622 580294 165678 580350
rect 165250 580170 165306 580226
rect 165374 580170 165430 580226
rect 165498 580170 165554 580226
rect 165622 580170 165678 580226
rect 165250 580046 165306 580102
rect 165374 580046 165430 580102
rect 165498 580046 165554 580102
rect 165622 580046 165678 580102
rect 165250 579922 165306 579978
rect 165374 579922 165430 579978
rect 165498 579922 165554 579978
rect 165622 579922 165678 579978
rect 165250 562294 165306 562350
rect 165374 562294 165430 562350
rect 165498 562294 165554 562350
rect 165622 562294 165678 562350
rect 165250 562170 165306 562226
rect 165374 562170 165430 562226
rect 165498 562170 165554 562226
rect 165622 562170 165678 562226
rect 165250 562046 165306 562102
rect 165374 562046 165430 562102
rect 165498 562046 165554 562102
rect 165622 562046 165678 562102
rect 165250 561922 165306 561978
rect 165374 561922 165430 561978
rect 165498 561922 165554 561978
rect 165622 561922 165678 561978
rect 165250 544294 165306 544350
rect 165374 544294 165430 544350
rect 165498 544294 165554 544350
rect 165622 544294 165678 544350
rect 165250 544170 165306 544226
rect 165374 544170 165430 544226
rect 165498 544170 165554 544226
rect 165622 544170 165678 544226
rect 165250 544046 165306 544102
rect 165374 544046 165430 544102
rect 165498 544046 165554 544102
rect 165622 544046 165678 544102
rect 165250 543922 165306 543978
rect 165374 543922 165430 543978
rect 165498 543922 165554 543978
rect 165622 543922 165678 543978
rect 165250 526294 165306 526350
rect 165374 526294 165430 526350
rect 165498 526294 165554 526350
rect 165622 526294 165678 526350
rect 165250 526170 165306 526226
rect 165374 526170 165430 526226
rect 165498 526170 165554 526226
rect 165622 526170 165678 526226
rect 165250 526046 165306 526102
rect 165374 526046 165430 526102
rect 165498 526046 165554 526102
rect 165622 526046 165678 526102
rect 165250 525922 165306 525978
rect 165374 525922 165430 525978
rect 165498 525922 165554 525978
rect 165622 525922 165678 525978
rect 168970 598116 169026 598172
rect 169094 598116 169150 598172
rect 169218 598116 169274 598172
rect 169342 598116 169398 598172
rect 168970 597992 169026 598048
rect 169094 597992 169150 598048
rect 169218 597992 169274 598048
rect 169342 597992 169398 598048
rect 168970 597868 169026 597924
rect 169094 597868 169150 597924
rect 169218 597868 169274 597924
rect 169342 597868 169398 597924
rect 168970 597744 169026 597800
rect 169094 597744 169150 597800
rect 169218 597744 169274 597800
rect 169342 597744 169398 597800
rect 168970 586294 169026 586350
rect 169094 586294 169150 586350
rect 169218 586294 169274 586350
rect 169342 586294 169398 586350
rect 168970 586170 169026 586226
rect 169094 586170 169150 586226
rect 169218 586170 169274 586226
rect 169342 586170 169398 586226
rect 168970 586046 169026 586102
rect 169094 586046 169150 586102
rect 169218 586046 169274 586102
rect 169342 586046 169398 586102
rect 168970 585922 169026 585978
rect 169094 585922 169150 585978
rect 169218 585922 169274 585978
rect 169342 585922 169398 585978
rect 168970 568294 169026 568350
rect 169094 568294 169150 568350
rect 169218 568294 169274 568350
rect 169342 568294 169398 568350
rect 168970 568170 169026 568226
rect 169094 568170 169150 568226
rect 169218 568170 169274 568226
rect 169342 568170 169398 568226
rect 168970 568046 169026 568102
rect 169094 568046 169150 568102
rect 169218 568046 169274 568102
rect 169342 568046 169398 568102
rect 168970 567922 169026 567978
rect 169094 567922 169150 567978
rect 169218 567922 169274 567978
rect 169342 567922 169398 567978
rect 168970 550294 169026 550350
rect 169094 550294 169150 550350
rect 169218 550294 169274 550350
rect 169342 550294 169398 550350
rect 168970 550170 169026 550226
rect 169094 550170 169150 550226
rect 169218 550170 169274 550226
rect 169342 550170 169398 550226
rect 168970 550046 169026 550102
rect 169094 550046 169150 550102
rect 169218 550046 169274 550102
rect 169342 550046 169398 550102
rect 168970 549922 169026 549978
rect 169094 549922 169150 549978
rect 169218 549922 169274 549978
rect 169342 549922 169398 549978
rect 168970 532294 169026 532350
rect 169094 532294 169150 532350
rect 169218 532294 169274 532350
rect 169342 532294 169398 532350
rect 168970 532170 169026 532226
rect 169094 532170 169150 532226
rect 169218 532170 169274 532226
rect 169342 532170 169398 532226
rect 168970 532046 169026 532102
rect 169094 532046 169150 532102
rect 169218 532046 169274 532102
rect 169342 532046 169398 532102
rect 168970 531922 169026 531978
rect 169094 531922 169150 531978
rect 169218 531922 169274 531978
rect 169342 531922 169398 531978
rect 183250 597156 183306 597212
rect 183374 597156 183430 597212
rect 183498 597156 183554 597212
rect 183622 597156 183678 597212
rect 183250 597032 183306 597088
rect 183374 597032 183430 597088
rect 183498 597032 183554 597088
rect 183622 597032 183678 597088
rect 183250 596908 183306 596964
rect 183374 596908 183430 596964
rect 183498 596908 183554 596964
rect 183622 596908 183678 596964
rect 183250 596784 183306 596840
rect 183374 596784 183430 596840
rect 183498 596784 183554 596840
rect 183622 596784 183678 596840
rect 183250 580294 183306 580350
rect 183374 580294 183430 580350
rect 183498 580294 183554 580350
rect 183622 580294 183678 580350
rect 183250 580170 183306 580226
rect 183374 580170 183430 580226
rect 183498 580170 183554 580226
rect 183622 580170 183678 580226
rect 183250 580046 183306 580102
rect 183374 580046 183430 580102
rect 183498 580046 183554 580102
rect 183622 580046 183678 580102
rect 183250 579922 183306 579978
rect 183374 579922 183430 579978
rect 183498 579922 183554 579978
rect 183622 579922 183678 579978
rect 183250 562294 183306 562350
rect 183374 562294 183430 562350
rect 183498 562294 183554 562350
rect 183622 562294 183678 562350
rect 183250 562170 183306 562226
rect 183374 562170 183430 562226
rect 183498 562170 183554 562226
rect 183622 562170 183678 562226
rect 183250 562046 183306 562102
rect 183374 562046 183430 562102
rect 183498 562046 183554 562102
rect 183622 562046 183678 562102
rect 183250 561922 183306 561978
rect 183374 561922 183430 561978
rect 183498 561922 183554 561978
rect 183622 561922 183678 561978
rect 183250 544294 183306 544350
rect 183374 544294 183430 544350
rect 183498 544294 183554 544350
rect 183622 544294 183678 544350
rect 183250 544170 183306 544226
rect 183374 544170 183430 544226
rect 183498 544170 183554 544226
rect 183622 544170 183678 544226
rect 183250 544046 183306 544102
rect 183374 544046 183430 544102
rect 183498 544046 183554 544102
rect 183622 544046 183678 544102
rect 183250 543922 183306 543978
rect 183374 543922 183430 543978
rect 183498 543922 183554 543978
rect 183622 543922 183678 543978
rect 183250 526294 183306 526350
rect 183374 526294 183430 526350
rect 183498 526294 183554 526350
rect 183622 526294 183678 526350
rect 183250 526170 183306 526226
rect 183374 526170 183430 526226
rect 183498 526170 183554 526226
rect 183622 526170 183678 526226
rect 183250 526046 183306 526102
rect 183374 526046 183430 526102
rect 183498 526046 183554 526102
rect 183622 526046 183678 526102
rect 183250 525922 183306 525978
rect 183374 525922 183430 525978
rect 183498 525922 183554 525978
rect 183622 525922 183678 525978
rect 186970 598116 187026 598172
rect 187094 598116 187150 598172
rect 187218 598116 187274 598172
rect 187342 598116 187398 598172
rect 186970 597992 187026 598048
rect 187094 597992 187150 598048
rect 187218 597992 187274 598048
rect 187342 597992 187398 598048
rect 186970 597868 187026 597924
rect 187094 597868 187150 597924
rect 187218 597868 187274 597924
rect 187342 597868 187398 597924
rect 186970 597744 187026 597800
rect 187094 597744 187150 597800
rect 187218 597744 187274 597800
rect 187342 597744 187398 597800
rect 186970 586294 187026 586350
rect 187094 586294 187150 586350
rect 187218 586294 187274 586350
rect 187342 586294 187398 586350
rect 186970 586170 187026 586226
rect 187094 586170 187150 586226
rect 187218 586170 187274 586226
rect 187342 586170 187398 586226
rect 186970 586046 187026 586102
rect 187094 586046 187150 586102
rect 187218 586046 187274 586102
rect 187342 586046 187398 586102
rect 186970 585922 187026 585978
rect 187094 585922 187150 585978
rect 187218 585922 187274 585978
rect 187342 585922 187398 585978
rect 186970 568294 187026 568350
rect 187094 568294 187150 568350
rect 187218 568294 187274 568350
rect 187342 568294 187398 568350
rect 186970 568170 187026 568226
rect 187094 568170 187150 568226
rect 187218 568170 187274 568226
rect 187342 568170 187398 568226
rect 186970 568046 187026 568102
rect 187094 568046 187150 568102
rect 187218 568046 187274 568102
rect 187342 568046 187398 568102
rect 186970 567922 187026 567978
rect 187094 567922 187150 567978
rect 187218 567922 187274 567978
rect 187342 567922 187398 567978
rect 186970 550294 187026 550350
rect 187094 550294 187150 550350
rect 187218 550294 187274 550350
rect 187342 550294 187398 550350
rect 186970 550170 187026 550226
rect 187094 550170 187150 550226
rect 187218 550170 187274 550226
rect 187342 550170 187398 550226
rect 186970 550046 187026 550102
rect 187094 550046 187150 550102
rect 187218 550046 187274 550102
rect 187342 550046 187398 550102
rect 186970 549922 187026 549978
rect 187094 549922 187150 549978
rect 187218 549922 187274 549978
rect 187342 549922 187398 549978
rect 186970 532294 187026 532350
rect 187094 532294 187150 532350
rect 187218 532294 187274 532350
rect 187342 532294 187398 532350
rect 186970 532170 187026 532226
rect 187094 532170 187150 532226
rect 187218 532170 187274 532226
rect 187342 532170 187398 532226
rect 186970 532046 187026 532102
rect 187094 532046 187150 532102
rect 187218 532046 187274 532102
rect 187342 532046 187398 532102
rect 186970 531922 187026 531978
rect 187094 531922 187150 531978
rect 187218 531922 187274 531978
rect 187342 531922 187398 531978
rect 201250 597156 201306 597212
rect 201374 597156 201430 597212
rect 201498 597156 201554 597212
rect 201622 597156 201678 597212
rect 201250 597032 201306 597088
rect 201374 597032 201430 597088
rect 201498 597032 201554 597088
rect 201622 597032 201678 597088
rect 201250 596908 201306 596964
rect 201374 596908 201430 596964
rect 201498 596908 201554 596964
rect 201622 596908 201678 596964
rect 201250 596784 201306 596840
rect 201374 596784 201430 596840
rect 201498 596784 201554 596840
rect 201622 596784 201678 596840
rect 201250 580294 201306 580350
rect 201374 580294 201430 580350
rect 201498 580294 201554 580350
rect 201622 580294 201678 580350
rect 201250 580170 201306 580226
rect 201374 580170 201430 580226
rect 201498 580170 201554 580226
rect 201622 580170 201678 580226
rect 201250 580046 201306 580102
rect 201374 580046 201430 580102
rect 201498 580046 201554 580102
rect 201622 580046 201678 580102
rect 201250 579922 201306 579978
rect 201374 579922 201430 579978
rect 201498 579922 201554 579978
rect 201622 579922 201678 579978
rect 201250 562294 201306 562350
rect 201374 562294 201430 562350
rect 201498 562294 201554 562350
rect 201622 562294 201678 562350
rect 201250 562170 201306 562226
rect 201374 562170 201430 562226
rect 201498 562170 201554 562226
rect 201622 562170 201678 562226
rect 201250 562046 201306 562102
rect 201374 562046 201430 562102
rect 201498 562046 201554 562102
rect 201622 562046 201678 562102
rect 201250 561922 201306 561978
rect 201374 561922 201430 561978
rect 201498 561922 201554 561978
rect 201622 561922 201678 561978
rect 201250 544294 201306 544350
rect 201374 544294 201430 544350
rect 201498 544294 201554 544350
rect 201622 544294 201678 544350
rect 201250 544170 201306 544226
rect 201374 544170 201430 544226
rect 201498 544170 201554 544226
rect 201622 544170 201678 544226
rect 201250 544046 201306 544102
rect 201374 544046 201430 544102
rect 201498 544046 201554 544102
rect 201622 544046 201678 544102
rect 201250 543922 201306 543978
rect 201374 543922 201430 543978
rect 201498 543922 201554 543978
rect 201622 543922 201678 543978
rect 201250 526294 201306 526350
rect 201374 526294 201430 526350
rect 201498 526294 201554 526350
rect 201622 526294 201678 526350
rect 201250 526170 201306 526226
rect 201374 526170 201430 526226
rect 201498 526170 201554 526226
rect 201622 526170 201678 526226
rect 201250 526046 201306 526102
rect 201374 526046 201430 526102
rect 201498 526046 201554 526102
rect 201622 526046 201678 526102
rect 201250 525922 201306 525978
rect 201374 525922 201430 525978
rect 201498 525922 201554 525978
rect 201622 525922 201678 525978
rect 204970 598116 205026 598172
rect 205094 598116 205150 598172
rect 205218 598116 205274 598172
rect 205342 598116 205398 598172
rect 204970 597992 205026 598048
rect 205094 597992 205150 598048
rect 205218 597992 205274 598048
rect 205342 597992 205398 598048
rect 204970 597868 205026 597924
rect 205094 597868 205150 597924
rect 205218 597868 205274 597924
rect 205342 597868 205398 597924
rect 204970 597744 205026 597800
rect 205094 597744 205150 597800
rect 205218 597744 205274 597800
rect 205342 597744 205398 597800
rect 204970 586294 205026 586350
rect 205094 586294 205150 586350
rect 205218 586294 205274 586350
rect 205342 586294 205398 586350
rect 204970 586170 205026 586226
rect 205094 586170 205150 586226
rect 205218 586170 205274 586226
rect 205342 586170 205398 586226
rect 204970 586046 205026 586102
rect 205094 586046 205150 586102
rect 205218 586046 205274 586102
rect 205342 586046 205398 586102
rect 204970 585922 205026 585978
rect 205094 585922 205150 585978
rect 205218 585922 205274 585978
rect 205342 585922 205398 585978
rect 204970 568294 205026 568350
rect 205094 568294 205150 568350
rect 205218 568294 205274 568350
rect 205342 568294 205398 568350
rect 204970 568170 205026 568226
rect 205094 568170 205150 568226
rect 205218 568170 205274 568226
rect 205342 568170 205398 568226
rect 204970 568046 205026 568102
rect 205094 568046 205150 568102
rect 205218 568046 205274 568102
rect 205342 568046 205398 568102
rect 204970 567922 205026 567978
rect 205094 567922 205150 567978
rect 205218 567922 205274 567978
rect 205342 567922 205398 567978
rect 204970 550294 205026 550350
rect 205094 550294 205150 550350
rect 205218 550294 205274 550350
rect 205342 550294 205398 550350
rect 204970 550170 205026 550226
rect 205094 550170 205150 550226
rect 205218 550170 205274 550226
rect 205342 550170 205398 550226
rect 204970 550046 205026 550102
rect 205094 550046 205150 550102
rect 205218 550046 205274 550102
rect 205342 550046 205398 550102
rect 204970 549922 205026 549978
rect 205094 549922 205150 549978
rect 205218 549922 205274 549978
rect 205342 549922 205398 549978
rect 204970 532294 205026 532350
rect 205094 532294 205150 532350
rect 205218 532294 205274 532350
rect 205342 532294 205398 532350
rect 204970 532170 205026 532226
rect 205094 532170 205150 532226
rect 205218 532170 205274 532226
rect 205342 532170 205398 532226
rect 204970 532046 205026 532102
rect 205094 532046 205150 532102
rect 205218 532046 205274 532102
rect 205342 532046 205398 532102
rect 204970 531922 205026 531978
rect 205094 531922 205150 531978
rect 205218 531922 205274 531978
rect 205342 531922 205398 531978
rect 219250 597156 219306 597212
rect 219374 597156 219430 597212
rect 219498 597156 219554 597212
rect 219622 597156 219678 597212
rect 219250 597032 219306 597088
rect 219374 597032 219430 597088
rect 219498 597032 219554 597088
rect 219622 597032 219678 597088
rect 219250 596908 219306 596964
rect 219374 596908 219430 596964
rect 219498 596908 219554 596964
rect 219622 596908 219678 596964
rect 219250 596784 219306 596840
rect 219374 596784 219430 596840
rect 219498 596784 219554 596840
rect 219622 596784 219678 596840
rect 219250 580294 219306 580350
rect 219374 580294 219430 580350
rect 219498 580294 219554 580350
rect 219622 580294 219678 580350
rect 219250 580170 219306 580226
rect 219374 580170 219430 580226
rect 219498 580170 219554 580226
rect 219622 580170 219678 580226
rect 219250 580046 219306 580102
rect 219374 580046 219430 580102
rect 219498 580046 219554 580102
rect 219622 580046 219678 580102
rect 219250 579922 219306 579978
rect 219374 579922 219430 579978
rect 219498 579922 219554 579978
rect 219622 579922 219678 579978
rect 219250 562294 219306 562350
rect 219374 562294 219430 562350
rect 219498 562294 219554 562350
rect 219622 562294 219678 562350
rect 219250 562170 219306 562226
rect 219374 562170 219430 562226
rect 219498 562170 219554 562226
rect 219622 562170 219678 562226
rect 219250 562046 219306 562102
rect 219374 562046 219430 562102
rect 219498 562046 219554 562102
rect 219622 562046 219678 562102
rect 219250 561922 219306 561978
rect 219374 561922 219430 561978
rect 219498 561922 219554 561978
rect 219622 561922 219678 561978
rect 219250 544294 219306 544350
rect 219374 544294 219430 544350
rect 219498 544294 219554 544350
rect 219622 544294 219678 544350
rect 219250 544170 219306 544226
rect 219374 544170 219430 544226
rect 219498 544170 219554 544226
rect 219622 544170 219678 544226
rect 219250 544046 219306 544102
rect 219374 544046 219430 544102
rect 219498 544046 219554 544102
rect 219622 544046 219678 544102
rect 219250 543922 219306 543978
rect 219374 543922 219430 543978
rect 219498 543922 219554 543978
rect 219622 543922 219678 543978
rect 219250 526294 219306 526350
rect 219374 526294 219430 526350
rect 219498 526294 219554 526350
rect 219622 526294 219678 526350
rect 219250 526170 219306 526226
rect 219374 526170 219430 526226
rect 219498 526170 219554 526226
rect 219622 526170 219678 526226
rect 219250 526046 219306 526102
rect 219374 526046 219430 526102
rect 219498 526046 219554 526102
rect 219622 526046 219678 526102
rect 219250 525922 219306 525978
rect 219374 525922 219430 525978
rect 219498 525922 219554 525978
rect 219622 525922 219678 525978
rect 222970 598116 223026 598172
rect 223094 598116 223150 598172
rect 223218 598116 223274 598172
rect 223342 598116 223398 598172
rect 222970 597992 223026 598048
rect 223094 597992 223150 598048
rect 223218 597992 223274 598048
rect 223342 597992 223398 598048
rect 222970 597868 223026 597924
rect 223094 597868 223150 597924
rect 223218 597868 223274 597924
rect 223342 597868 223398 597924
rect 222970 597744 223026 597800
rect 223094 597744 223150 597800
rect 223218 597744 223274 597800
rect 223342 597744 223398 597800
rect 222970 586294 223026 586350
rect 223094 586294 223150 586350
rect 223218 586294 223274 586350
rect 223342 586294 223398 586350
rect 222970 586170 223026 586226
rect 223094 586170 223150 586226
rect 223218 586170 223274 586226
rect 223342 586170 223398 586226
rect 222970 586046 223026 586102
rect 223094 586046 223150 586102
rect 223218 586046 223274 586102
rect 223342 586046 223398 586102
rect 222970 585922 223026 585978
rect 223094 585922 223150 585978
rect 223218 585922 223274 585978
rect 223342 585922 223398 585978
rect 222970 568294 223026 568350
rect 223094 568294 223150 568350
rect 223218 568294 223274 568350
rect 223342 568294 223398 568350
rect 222970 568170 223026 568226
rect 223094 568170 223150 568226
rect 223218 568170 223274 568226
rect 223342 568170 223398 568226
rect 222970 568046 223026 568102
rect 223094 568046 223150 568102
rect 223218 568046 223274 568102
rect 223342 568046 223398 568102
rect 222970 567922 223026 567978
rect 223094 567922 223150 567978
rect 223218 567922 223274 567978
rect 223342 567922 223398 567978
rect 222970 550294 223026 550350
rect 223094 550294 223150 550350
rect 223218 550294 223274 550350
rect 223342 550294 223398 550350
rect 222970 550170 223026 550226
rect 223094 550170 223150 550226
rect 223218 550170 223274 550226
rect 223342 550170 223398 550226
rect 222970 550046 223026 550102
rect 223094 550046 223150 550102
rect 223218 550046 223274 550102
rect 223342 550046 223398 550102
rect 222970 549922 223026 549978
rect 223094 549922 223150 549978
rect 223218 549922 223274 549978
rect 223342 549922 223398 549978
rect 222970 532294 223026 532350
rect 223094 532294 223150 532350
rect 223218 532294 223274 532350
rect 223342 532294 223398 532350
rect 222970 532170 223026 532226
rect 223094 532170 223150 532226
rect 223218 532170 223274 532226
rect 223342 532170 223398 532226
rect 222970 532046 223026 532102
rect 223094 532046 223150 532102
rect 223218 532046 223274 532102
rect 223342 532046 223398 532102
rect 222970 531922 223026 531978
rect 223094 531922 223150 531978
rect 223218 531922 223274 531978
rect 223342 531922 223398 531978
rect 237250 597156 237306 597212
rect 237374 597156 237430 597212
rect 237498 597156 237554 597212
rect 237622 597156 237678 597212
rect 237250 597032 237306 597088
rect 237374 597032 237430 597088
rect 237498 597032 237554 597088
rect 237622 597032 237678 597088
rect 237250 596908 237306 596964
rect 237374 596908 237430 596964
rect 237498 596908 237554 596964
rect 237622 596908 237678 596964
rect 237250 596784 237306 596840
rect 237374 596784 237430 596840
rect 237498 596784 237554 596840
rect 237622 596784 237678 596840
rect 237250 580294 237306 580350
rect 237374 580294 237430 580350
rect 237498 580294 237554 580350
rect 237622 580294 237678 580350
rect 237250 580170 237306 580226
rect 237374 580170 237430 580226
rect 237498 580170 237554 580226
rect 237622 580170 237678 580226
rect 237250 580046 237306 580102
rect 237374 580046 237430 580102
rect 237498 580046 237554 580102
rect 237622 580046 237678 580102
rect 237250 579922 237306 579978
rect 237374 579922 237430 579978
rect 237498 579922 237554 579978
rect 237622 579922 237678 579978
rect 237250 562294 237306 562350
rect 237374 562294 237430 562350
rect 237498 562294 237554 562350
rect 237622 562294 237678 562350
rect 237250 562170 237306 562226
rect 237374 562170 237430 562226
rect 237498 562170 237554 562226
rect 237622 562170 237678 562226
rect 237250 562046 237306 562102
rect 237374 562046 237430 562102
rect 237498 562046 237554 562102
rect 237622 562046 237678 562102
rect 237250 561922 237306 561978
rect 237374 561922 237430 561978
rect 237498 561922 237554 561978
rect 237622 561922 237678 561978
rect 237250 544294 237306 544350
rect 237374 544294 237430 544350
rect 237498 544294 237554 544350
rect 237622 544294 237678 544350
rect 237250 544170 237306 544226
rect 237374 544170 237430 544226
rect 237498 544170 237554 544226
rect 237622 544170 237678 544226
rect 237250 544046 237306 544102
rect 237374 544046 237430 544102
rect 237498 544046 237554 544102
rect 237622 544046 237678 544102
rect 237250 543922 237306 543978
rect 237374 543922 237430 543978
rect 237498 543922 237554 543978
rect 237622 543922 237678 543978
rect 237250 526294 237306 526350
rect 237374 526294 237430 526350
rect 237498 526294 237554 526350
rect 237622 526294 237678 526350
rect 237250 526170 237306 526226
rect 237374 526170 237430 526226
rect 237498 526170 237554 526226
rect 237622 526170 237678 526226
rect 237250 526046 237306 526102
rect 237374 526046 237430 526102
rect 237498 526046 237554 526102
rect 237622 526046 237678 526102
rect 237250 525922 237306 525978
rect 237374 525922 237430 525978
rect 237498 525922 237554 525978
rect 237622 525922 237678 525978
rect 240970 598116 241026 598172
rect 241094 598116 241150 598172
rect 241218 598116 241274 598172
rect 241342 598116 241398 598172
rect 240970 597992 241026 598048
rect 241094 597992 241150 598048
rect 241218 597992 241274 598048
rect 241342 597992 241398 598048
rect 240970 597868 241026 597924
rect 241094 597868 241150 597924
rect 241218 597868 241274 597924
rect 241342 597868 241398 597924
rect 240970 597744 241026 597800
rect 241094 597744 241150 597800
rect 241218 597744 241274 597800
rect 241342 597744 241398 597800
rect 240970 586294 241026 586350
rect 241094 586294 241150 586350
rect 241218 586294 241274 586350
rect 241342 586294 241398 586350
rect 240970 586170 241026 586226
rect 241094 586170 241150 586226
rect 241218 586170 241274 586226
rect 241342 586170 241398 586226
rect 240970 586046 241026 586102
rect 241094 586046 241150 586102
rect 241218 586046 241274 586102
rect 241342 586046 241398 586102
rect 240970 585922 241026 585978
rect 241094 585922 241150 585978
rect 241218 585922 241274 585978
rect 241342 585922 241398 585978
rect 240970 568294 241026 568350
rect 241094 568294 241150 568350
rect 241218 568294 241274 568350
rect 241342 568294 241398 568350
rect 240970 568170 241026 568226
rect 241094 568170 241150 568226
rect 241218 568170 241274 568226
rect 241342 568170 241398 568226
rect 240970 568046 241026 568102
rect 241094 568046 241150 568102
rect 241218 568046 241274 568102
rect 241342 568046 241398 568102
rect 240970 567922 241026 567978
rect 241094 567922 241150 567978
rect 241218 567922 241274 567978
rect 241342 567922 241398 567978
rect 240970 550294 241026 550350
rect 241094 550294 241150 550350
rect 241218 550294 241274 550350
rect 241342 550294 241398 550350
rect 240970 550170 241026 550226
rect 241094 550170 241150 550226
rect 241218 550170 241274 550226
rect 241342 550170 241398 550226
rect 240970 550046 241026 550102
rect 241094 550046 241150 550102
rect 241218 550046 241274 550102
rect 241342 550046 241398 550102
rect 240970 549922 241026 549978
rect 241094 549922 241150 549978
rect 241218 549922 241274 549978
rect 241342 549922 241398 549978
rect 240970 532294 241026 532350
rect 241094 532294 241150 532350
rect 241218 532294 241274 532350
rect 241342 532294 241398 532350
rect 240970 532170 241026 532226
rect 241094 532170 241150 532226
rect 241218 532170 241274 532226
rect 241342 532170 241398 532226
rect 240970 532046 241026 532102
rect 241094 532046 241150 532102
rect 241218 532046 241274 532102
rect 241342 532046 241398 532102
rect 240970 531922 241026 531978
rect 241094 531922 241150 531978
rect 241218 531922 241274 531978
rect 241342 531922 241398 531978
rect 255250 597156 255306 597212
rect 255374 597156 255430 597212
rect 255498 597156 255554 597212
rect 255622 597156 255678 597212
rect 255250 597032 255306 597088
rect 255374 597032 255430 597088
rect 255498 597032 255554 597088
rect 255622 597032 255678 597088
rect 255250 596908 255306 596964
rect 255374 596908 255430 596964
rect 255498 596908 255554 596964
rect 255622 596908 255678 596964
rect 255250 596784 255306 596840
rect 255374 596784 255430 596840
rect 255498 596784 255554 596840
rect 255622 596784 255678 596840
rect 255250 580294 255306 580350
rect 255374 580294 255430 580350
rect 255498 580294 255554 580350
rect 255622 580294 255678 580350
rect 255250 580170 255306 580226
rect 255374 580170 255430 580226
rect 255498 580170 255554 580226
rect 255622 580170 255678 580226
rect 255250 580046 255306 580102
rect 255374 580046 255430 580102
rect 255498 580046 255554 580102
rect 255622 580046 255678 580102
rect 255250 579922 255306 579978
rect 255374 579922 255430 579978
rect 255498 579922 255554 579978
rect 255622 579922 255678 579978
rect 255250 562294 255306 562350
rect 255374 562294 255430 562350
rect 255498 562294 255554 562350
rect 255622 562294 255678 562350
rect 255250 562170 255306 562226
rect 255374 562170 255430 562226
rect 255498 562170 255554 562226
rect 255622 562170 255678 562226
rect 255250 562046 255306 562102
rect 255374 562046 255430 562102
rect 255498 562046 255554 562102
rect 255622 562046 255678 562102
rect 255250 561922 255306 561978
rect 255374 561922 255430 561978
rect 255498 561922 255554 561978
rect 255622 561922 255678 561978
rect 255250 544294 255306 544350
rect 255374 544294 255430 544350
rect 255498 544294 255554 544350
rect 255622 544294 255678 544350
rect 255250 544170 255306 544226
rect 255374 544170 255430 544226
rect 255498 544170 255554 544226
rect 255622 544170 255678 544226
rect 255250 544046 255306 544102
rect 255374 544046 255430 544102
rect 255498 544046 255554 544102
rect 255622 544046 255678 544102
rect 255250 543922 255306 543978
rect 255374 543922 255430 543978
rect 255498 543922 255554 543978
rect 255622 543922 255678 543978
rect 255250 526294 255306 526350
rect 255374 526294 255430 526350
rect 255498 526294 255554 526350
rect 255622 526294 255678 526350
rect 255250 526170 255306 526226
rect 255374 526170 255430 526226
rect 255498 526170 255554 526226
rect 255622 526170 255678 526226
rect 255250 526046 255306 526102
rect 255374 526046 255430 526102
rect 255498 526046 255554 526102
rect 255622 526046 255678 526102
rect 255250 525922 255306 525978
rect 255374 525922 255430 525978
rect 255498 525922 255554 525978
rect 255622 525922 255678 525978
rect 258970 598116 259026 598172
rect 259094 598116 259150 598172
rect 259218 598116 259274 598172
rect 259342 598116 259398 598172
rect 258970 597992 259026 598048
rect 259094 597992 259150 598048
rect 259218 597992 259274 598048
rect 259342 597992 259398 598048
rect 258970 597868 259026 597924
rect 259094 597868 259150 597924
rect 259218 597868 259274 597924
rect 259342 597868 259398 597924
rect 258970 597744 259026 597800
rect 259094 597744 259150 597800
rect 259218 597744 259274 597800
rect 259342 597744 259398 597800
rect 258970 586294 259026 586350
rect 259094 586294 259150 586350
rect 259218 586294 259274 586350
rect 259342 586294 259398 586350
rect 258970 586170 259026 586226
rect 259094 586170 259150 586226
rect 259218 586170 259274 586226
rect 259342 586170 259398 586226
rect 258970 586046 259026 586102
rect 259094 586046 259150 586102
rect 259218 586046 259274 586102
rect 259342 586046 259398 586102
rect 258970 585922 259026 585978
rect 259094 585922 259150 585978
rect 259218 585922 259274 585978
rect 259342 585922 259398 585978
rect 258970 568294 259026 568350
rect 259094 568294 259150 568350
rect 259218 568294 259274 568350
rect 259342 568294 259398 568350
rect 258970 568170 259026 568226
rect 259094 568170 259150 568226
rect 259218 568170 259274 568226
rect 259342 568170 259398 568226
rect 258970 568046 259026 568102
rect 259094 568046 259150 568102
rect 259218 568046 259274 568102
rect 259342 568046 259398 568102
rect 258970 567922 259026 567978
rect 259094 567922 259150 567978
rect 259218 567922 259274 567978
rect 259342 567922 259398 567978
rect 258970 550294 259026 550350
rect 259094 550294 259150 550350
rect 259218 550294 259274 550350
rect 259342 550294 259398 550350
rect 258970 550170 259026 550226
rect 259094 550170 259150 550226
rect 259218 550170 259274 550226
rect 259342 550170 259398 550226
rect 258970 550046 259026 550102
rect 259094 550046 259150 550102
rect 259218 550046 259274 550102
rect 259342 550046 259398 550102
rect 258970 549922 259026 549978
rect 259094 549922 259150 549978
rect 259218 549922 259274 549978
rect 259342 549922 259398 549978
rect 258970 532294 259026 532350
rect 259094 532294 259150 532350
rect 259218 532294 259274 532350
rect 259342 532294 259398 532350
rect 258970 532170 259026 532226
rect 259094 532170 259150 532226
rect 259218 532170 259274 532226
rect 259342 532170 259398 532226
rect 258970 532046 259026 532102
rect 259094 532046 259150 532102
rect 259218 532046 259274 532102
rect 259342 532046 259398 532102
rect 258970 531922 259026 531978
rect 259094 531922 259150 531978
rect 259218 531922 259274 531978
rect 259342 531922 259398 531978
rect 273250 597156 273306 597212
rect 273374 597156 273430 597212
rect 273498 597156 273554 597212
rect 273622 597156 273678 597212
rect 273250 597032 273306 597088
rect 273374 597032 273430 597088
rect 273498 597032 273554 597088
rect 273622 597032 273678 597088
rect 273250 596908 273306 596964
rect 273374 596908 273430 596964
rect 273498 596908 273554 596964
rect 273622 596908 273678 596964
rect 273250 596784 273306 596840
rect 273374 596784 273430 596840
rect 273498 596784 273554 596840
rect 273622 596784 273678 596840
rect 273250 580294 273306 580350
rect 273374 580294 273430 580350
rect 273498 580294 273554 580350
rect 273622 580294 273678 580350
rect 273250 580170 273306 580226
rect 273374 580170 273430 580226
rect 273498 580170 273554 580226
rect 273622 580170 273678 580226
rect 273250 580046 273306 580102
rect 273374 580046 273430 580102
rect 273498 580046 273554 580102
rect 273622 580046 273678 580102
rect 273250 579922 273306 579978
rect 273374 579922 273430 579978
rect 273498 579922 273554 579978
rect 273622 579922 273678 579978
rect 273250 562294 273306 562350
rect 273374 562294 273430 562350
rect 273498 562294 273554 562350
rect 273622 562294 273678 562350
rect 273250 562170 273306 562226
rect 273374 562170 273430 562226
rect 273498 562170 273554 562226
rect 273622 562170 273678 562226
rect 273250 562046 273306 562102
rect 273374 562046 273430 562102
rect 273498 562046 273554 562102
rect 273622 562046 273678 562102
rect 273250 561922 273306 561978
rect 273374 561922 273430 561978
rect 273498 561922 273554 561978
rect 273622 561922 273678 561978
rect 273250 544294 273306 544350
rect 273374 544294 273430 544350
rect 273498 544294 273554 544350
rect 273622 544294 273678 544350
rect 273250 544170 273306 544226
rect 273374 544170 273430 544226
rect 273498 544170 273554 544226
rect 273622 544170 273678 544226
rect 273250 544046 273306 544102
rect 273374 544046 273430 544102
rect 273498 544046 273554 544102
rect 273622 544046 273678 544102
rect 273250 543922 273306 543978
rect 273374 543922 273430 543978
rect 273498 543922 273554 543978
rect 273622 543922 273678 543978
rect 273250 526294 273306 526350
rect 273374 526294 273430 526350
rect 273498 526294 273554 526350
rect 273622 526294 273678 526350
rect 273250 526170 273306 526226
rect 273374 526170 273430 526226
rect 273498 526170 273554 526226
rect 273622 526170 273678 526226
rect 273250 526046 273306 526102
rect 273374 526046 273430 526102
rect 273498 526046 273554 526102
rect 273622 526046 273678 526102
rect 273250 525922 273306 525978
rect 273374 525922 273430 525978
rect 273498 525922 273554 525978
rect 273622 525922 273678 525978
rect 276970 598116 277026 598172
rect 277094 598116 277150 598172
rect 277218 598116 277274 598172
rect 277342 598116 277398 598172
rect 276970 597992 277026 598048
rect 277094 597992 277150 598048
rect 277218 597992 277274 598048
rect 277342 597992 277398 598048
rect 276970 597868 277026 597924
rect 277094 597868 277150 597924
rect 277218 597868 277274 597924
rect 277342 597868 277398 597924
rect 276970 597744 277026 597800
rect 277094 597744 277150 597800
rect 277218 597744 277274 597800
rect 277342 597744 277398 597800
rect 276970 586294 277026 586350
rect 277094 586294 277150 586350
rect 277218 586294 277274 586350
rect 277342 586294 277398 586350
rect 276970 586170 277026 586226
rect 277094 586170 277150 586226
rect 277218 586170 277274 586226
rect 277342 586170 277398 586226
rect 276970 586046 277026 586102
rect 277094 586046 277150 586102
rect 277218 586046 277274 586102
rect 277342 586046 277398 586102
rect 276970 585922 277026 585978
rect 277094 585922 277150 585978
rect 277218 585922 277274 585978
rect 277342 585922 277398 585978
rect 276970 568294 277026 568350
rect 277094 568294 277150 568350
rect 277218 568294 277274 568350
rect 277342 568294 277398 568350
rect 276970 568170 277026 568226
rect 277094 568170 277150 568226
rect 277218 568170 277274 568226
rect 277342 568170 277398 568226
rect 276970 568046 277026 568102
rect 277094 568046 277150 568102
rect 277218 568046 277274 568102
rect 277342 568046 277398 568102
rect 276970 567922 277026 567978
rect 277094 567922 277150 567978
rect 277218 567922 277274 567978
rect 277342 567922 277398 567978
rect 276970 550294 277026 550350
rect 277094 550294 277150 550350
rect 277218 550294 277274 550350
rect 277342 550294 277398 550350
rect 276970 550170 277026 550226
rect 277094 550170 277150 550226
rect 277218 550170 277274 550226
rect 277342 550170 277398 550226
rect 276970 550046 277026 550102
rect 277094 550046 277150 550102
rect 277218 550046 277274 550102
rect 277342 550046 277398 550102
rect 276970 549922 277026 549978
rect 277094 549922 277150 549978
rect 277218 549922 277274 549978
rect 277342 549922 277398 549978
rect 276970 532294 277026 532350
rect 277094 532294 277150 532350
rect 277218 532294 277274 532350
rect 277342 532294 277398 532350
rect 276970 532170 277026 532226
rect 277094 532170 277150 532226
rect 277218 532170 277274 532226
rect 277342 532170 277398 532226
rect 276970 532046 277026 532102
rect 277094 532046 277150 532102
rect 277218 532046 277274 532102
rect 277342 532046 277398 532102
rect 276970 531922 277026 531978
rect 277094 531922 277150 531978
rect 277218 531922 277274 531978
rect 277342 531922 277398 531978
rect 291250 597156 291306 597212
rect 291374 597156 291430 597212
rect 291498 597156 291554 597212
rect 291622 597156 291678 597212
rect 291250 597032 291306 597088
rect 291374 597032 291430 597088
rect 291498 597032 291554 597088
rect 291622 597032 291678 597088
rect 291250 596908 291306 596964
rect 291374 596908 291430 596964
rect 291498 596908 291554 596964
rect 291622 596908 291678 596964
rect 291250 596784 291306 596840
rect 291374 596784 291430 596840
rect 291498 596784 291554 596840
rect 291622 596784 291678 596840
rect 291250 580294 291306 580350
rect 291374 580294 291430 580350
rect 291498 580294 291554 580350
rect 291622 580294 291678 580350
rect 291250 580170 291306 580226
rect 291374 580170 291430 580226
rect 291498 580170 291554 580226
rect 291622 580170 291678 580226
rect 291250 580046 291306 580102
rect 291374 580046 291430 580102
rect 291498 580046 291554 580102
rect 291622 580046 291678 580102
rect 291250 579922 291306 579978
rect 291374 579922 291430 579978
rect 291498 579922 291554 579978
rect 291622 579922 291678 579978
rect 291250 562294 291306 562350
rect 291374 562294 291430 562350
rect 291498 562294 291554 562350
rect 291622 562294 291678 562350
rect 291250 562170 291306 562226
rect 291374 562170 291430 562226
rect 291498 562170 291554 562226
rect 291622 562170 291678 562226
rect 291250 562046 291306 562102
rect 291374 562046 291430 562102
rect 291498 562046 291554 562102
rect 291622 562046 291678 562102
rect 291250 561922 291306 561978
rect 291374 561922 291430 561978
rect 291498 561922 291554 561978
rect 291622 561922 291678 561978
rect 291250 544294 291306 544350
rect 291374 544294 291430 544350
rect 291498 544294 291554 544350
rect 291622 544294 291678 544350
rect 291250 544170 291306 544226
rect 291374 544170 291430 544226
rect 291498 544170 291554 544226
rect 291622 544170 291678 544226
rect 291250 544046 291306 544102
rect 291374 544046 291430 544102
rect 291498 544046 291554 544102
rect 291622 544046 291678 544102
rect 291250 543922 291306 543978
rect 291374 543922 291430 543978
rect 291498 543922 291554 543978
rect 291622 543922 291678 543978
rect 291250 526294 291306 526350
rect 291374 526294 291430 526350
rect 291498 526294 291554 526350
rect 291622 526294 291678 526350
rect 291250 526170 291306 526226
rect 291374 526170 291430 526226
rect 291498 526170 291554 526226
rect 291622 526170 291678 526226
rect 291250 526046 291306 526102
rect 291374 526046 291430 526102
rect 291498 526046 291554 526102
rect 291622 526046 291678 526102
rect 291250 525922 291306 525978
rect 291374 525922 291430 525978
rect 291498 525922 291554 525978
rect 291622 525922 291678 525978
rect 294970 598116 295026 598172
rect 295094 598116 295150 598172
rect 295218 598116 295274 598172
rect 295342 598116 295398 598172
rect 294970 597992 295026 598048
rect 295094 597992 295150 598048
rect 295218 597992 295274 598048
rect 295342 597992 295398 598048
rect 294970 597868 295026 597924
rect 295094 597868 295150 597924
rect 295218 597868 295274 597924
rect 295342 597868 295398 597924
rect 294970 597744 295026 597800
rect 295094 597744 295150 597800
rect 295218 597744 295274 597800
rect 295342 597744 295398 597800
rect 294970 586294 295026 586350
rect 295094 586294 295150 586350
rect 295218 586294 295274 586350
rect 295342 586294 295398 586350
rect 294970 586170 295026 586226
rect 295094 586170 295150 586226
rect 295218 586170 295274 586226
rect 295342 586170 295398 586226
rect 294970 586046 295026 586102
rect 295094 586046 295150 586102
rect 295218 586046 295274 586102
rect 295342 586046 295398 586102
rect 294970 585922 295026 585978
rect 295094 585922 295150 585978
rect 295218 585922 295274 585978
rect 295342 585922 295398 585978
rect 294970 568294 295026 568350
rect 295094 568294 295150 568350
rect 295218 568294 295274 568350
rect 295342 568294 295398 568350
rect 294970 568170 295026 568226
rect 295094 568170 295150 568226
rect 295218 568170 295274 568226
rect 295342 568170 295398 568226
rect 294970 568046 295026 568102
rect 295094 568046 295150 568102
rect 295218 568046 295274 568102
rect 295342 568046 295398 568102
rect 294970 567922 295026 567978
rect 295094 567922 295150 567978
rect 295218 567922 295274 567978
rect 295342 567922 295398 567978
rect 294970 550294 295026 550350
rect 295094 550294 295150 550350
rect 295218 550294 295274 550350
rect 295342 550294 295398 550350
rect 294970 550170 295026 550226
rect 295094 550170 295150 550226
rect 295218 550170 295274 550226
rect 295342 550170 295398 550226
rect 294970 550046 295026 550102
rect 295094 550046 295150 550102
rect 295218 550046 295274 550102
rect 295342 550046 295398 550102
rect 294970 549922 295026 549978
rect 295094 549922 295150 549978
rect 295218 549922 295274 549978
rect 295342 549922 295398 549978
rect 294970 532294 295026 532350
rect 295094 532294 295150 532350
rect 295218 532294 295274 532350
rect 295342 532294 295398 532350
rect 294970 532170 295026 532226
rect 295094 532170 295150 532226
rect 295218 532170 295274 532226
rect 295342 532170 295398 532226
rect 294970 532046 295026 532102
rect 295094 532046 295150 532102
rect 295218 532046 295274 532102
rect 295342 532046 295398 532102
rect 294970 531922 295026 531978
rect 295094 531922 295150 531978
rect 295218 531922 295274 531978
rect 295342 531922 295398 531978
rect 309250 597156 309306 597212
rect 309374 597156 309430 597212
rect 309498 597156 309554 597212
rect 309622 597156 309678 597212
rect 309250 597032 309306 597088
rect 309374 597032 309430 597088
rect 309498 597032 309554 597088
rect 309622 597032 309678 597088
rect 309250 596908 309306 596964
rect 309374 596908 309430 596964
rect 309498 596908 309554 596964
rect 309622 596908 309678 596964
rect 309250 596784 309306 596840
rect 309374 596784 309430 596840
rect 309498 596784 309554 596840
rect 309622 596784 309678 596840
rect 309250 580294 309306 580350
rect 309374 580294 309430 580350
rect 309498 580294 309554 580350
rect 309622 580294 309678 580350
rect 309250 580170 309306 580226
rect 309374 580170 309430 580226
rect 309498 580170 309554 580226
rect 309622 580170 309678 580226
rect 309250 580046 309306 580102
rect 309374 580046 309430 580102
rect 309498 580046 309554 580102
rect 309622 580046 309678 580102
rect 309250 579922 309306 579978
rect 309374 579922 309430 579978
rect 309498 579922 309554 579978
rect 309622 579922 309678 579978
rect 309250 562294 309306 562350
rect 309374 562294 309430 562350
rect 309498 562294 309554 562350
rect 309622 562294 309678 562350
rect 309250 562170 309306 562226
rect 309374 562170 309430 562226
rect 309498 562170 309554 562226
rect 309622 562170 309678 562226
rect 309250 562046 309306 562102
rect 309374 562046 309430 562102
rect 309498 562046 309554 562102
rect 309622 562046 309678 562102
rect 309250 561922 309306 561978
rect 309374 561922 309430 561978
rect 309498 561922 309554 561978
rect 309622 561922 309678 561978
rect 309250 544294 309306 544350
rect 309374 544294 309430 544350
rect 309498 544294 309554 544350
rect 309622 544294 309678 544350
rect 309250 544170 309306 544226
rect 309374 544170 309430 544226
rect 309498 544170 309554 544226
rect 309622 544170 309678 544226
rect 309250 544046 309306 544102
rect 309374 544046 309430 544102
rect 309498 544046 309554 544102
rect 309622 544046 309678 544102
rect 309250 543922 309306 543978
rect 309374 543922 309430 543978
rect 309498 543922 309554 543978
rect 309622 543922 309678 543978
rect 309250 526294 309306 526350
rect 309374 526294 309430 526350
rect 309498 526294 309554 526350
rect 309622 526294 309678 526350
rect 309250 526170 309306 526226
rect 309374 526170 309430 526226
rect 309498 526170 309554 526226
rect 309622 526170 309678 526226
rect 309250 526046 309306 526102
rect 309374 526046 309430 526102
rect 309498 526046 309554 526102
rect 309622 526046 309678 526102
rect 309250 525922 309306 525978
rect 309374 525922 309430 525978
rect 309498 525922 309554 525978
rect 309622 525922 309678 525978
rect 312970 598116 313026 598172
rect 313094 598116 313150 598172
rect 313218 598116 313274 598172
rect 313342 598116 313398 598172
rect 312970 597992 313026 598048
rect 313094 597992 313150 598048
rect 313218 597992 313274 598048
rect 313342 597992 313398 598048
rect 312970 597868 313026 597924
rect 313094 597868 313150 597924
rect 313218 597868 313274 597924
rect 313342 597868 313398 597924
rect 312970 597744 313026 597800
rect 313094 597744 313150 597800
rect 313218 597744 313274 597800
rect 313342 597744 313398 597800
rect 312970 586294 313026 586350
rect 313094 586294 313150 586350
rect 313218 586294 313274 586350
rect 313342 586294 313398 586350
rect 312970 586170 313026 586226
rect 313094 586170 313150 586226
rect 313218 586170 313274 586226
rect 313342 586170 313398 586226
rect 312970 586046 313026 586102
rect 313094 586046 313150 586102
rect 313218 586046 313274 586102
rect 313342 586046 313398 586102
rect 312970 585922 313026 585978
rect 313094 585922 313150 585978
rect 313218 585922 313274 585978
rect 313342 585922 313398 585978
rect 312970 568294 313026 568350
rect 313094 568294 313150 568350
rect 313218 568294 313274 568350
rect 313342 568294 313398 568350
rect 312970 568170 313026 568226
rect 313094 568170 313150 568226
rect 313218 568170 313274 568226
rect 313342 568170 313398 568226
rect 312970 568046 313026 568102
rect 313094 568046 313150 568102
rect 313218 568046 313274 568102
rect 313342 568046 313398 568102
rect 312970 567922 313026 567978
rect 313094 567922 313150 567978
rect 313218 567922 313274 567978
rect 313342 567922 313398 567978
rect 312970 550294 313026 550350
rect 313094 550294 313150 550350
rect 313218 550294 313274 550350
rect 313342 550294 313398 550350
rect 312970 550170 313026 550226
rect 313094 550170 313150 550226
rect 313218 550170 313274 550226
rect 313342 550170 313398 550226
rect 312970 550046 313026 550102
rect 313094 550046 313150 550102
rect 313218 550046 313274 550102
rect 313342 550046 313398 550102
rect 312970 549922 313026 549978
rect 313094 549922 313150 549978
rect 313218 549922 313274 549978
rect 313342 549922 313398 549978
rect 312970 532294 313026 532350
rect 313094 532294 313150 532350
rect 313218 532294 313274 532350
rect 313342 532294 313398 532350
rect 312970 532170 313026 532226
rect 313094 532170 313150 532226
rect 313218 532170 313274 532226
rect 313342 532170 313398 532226
rect 312970 532046 313026 532102
rect 313094 532046 313150 532102
rect 313218 532046 313274 532102
rect 313342 532046 313398 532102
rect 312970 531922 313026 531978
rect 313094 531922 313150 531978
rect 313218 531922 313274 531978
rect 313342 531922 313398 531978
rect 327250 597156 327306 597212
rect 327374 597156 327430 597212
rect 327498 597156 327554 597212
rect 327622 597156 327678 597212
rect 327250 597032 327306 597088
rect 327374 597032 327430 597088
rect 327498 597032 327554 597088
rect 327622 597032 327678 597088
rect 327250 596908 327306 596964
rect 327374 596908 327430 596964
rect 327498 596908 327554 596964
rect 327622 596908 327678 596964
rect 327250 596784 327306 596840
rect 327374 596784 327430 596840
rect 327498 596784 327554 596840
rect 327622 596784 327678 596840
rect 327250 580294 327306 580350
rect 327374 580294 327430 580350
rect 327498 580294 327554 580350
rect 327622 580294 327678 580350
rect 327250 580170 327306 580226
rect 327374 580170 327430 580226
rect 327498 580170 327554 580226
rect 327622 580170 327678 580226
rect 327250 580046 327306 580102
rect 327374 580046 327430 580102
rect 327498 580046 327554 580102
rect 327622 580046 327678 580102
rect 327250 579922 327306 579978
rect 327374 579922 327430 579978
rect 327498 579922 327554 579978
rect 327622 579922 327678 579978
rect 327250 562294 327306 562350
rect 327374 562294 327430 562350
rect 327498 562294 327554 562350
rect 327622 562294 327678 562350
rect 327250 562170 327306 562226
rect 327374 562170 327430 562226
rect 327498 562170 327554 562226
rect 327622 562170 327678 562226
rect 327250 562046 327306 562102
rect 327374 562046 327430 562102
rect 327498 562046 327554 562102
rect 327622 562046 327678 562102
rect 327250 561922 327306 561978
rect 327374 561922 327430 561978
rect 327498 561922 327554 561978
rect 327622 561922 327678 561978
rect 327250 544294 327306 544350
rect 327374 544294 327430 544350
rect 327498 544294 327554 544350
rect 327622 544294 327678 544350
rect 327250 544170 327306 544226
rect 327374 544170 327430 544226
rect 327498 544170 327554 544226
rect 327622 544170 327678 544226
rect 327250 544046 327306 544102
rect 327374 544046 327430 544102
rect 327498 544046 327554 544102
rect 327622 544046 327678 544102
rect 327250 543922 327306 543978
rect 327374 543922 327430 543978
rect 327498 543922 327554 543978
rect 327622 543922 327678 543978
rect 327250 526294 327306 526350
rect 327374 526294 327430 526350
rect 327498 526294 327554 526350
rect 327622 526294 327678 526350
rect 327250 526170 327306 526226
rect 327374 526170 327430 526226
rect 327498 526170 327554 526226
rect 327622 526170 327678 526226
rect 327250 526046 327306 526102
rect 327374 526046 327430 526102
rect 327498 526046 327554 526102
rect 327622 526046 327678 526102
rect 327250 525922 327306 525978
rect 327374 525922 327430 525978
rect 327498 525922 327554 525978
rect 327622 525922 327678 525978
rect 330970 598116 331026 598172
rect 331094 598116 331150 598172
rect 331218 598116 331274 598172
rect 331342 598116 331398 598172
rect 330970 597992 331026 598048
rect 331094 597992 331150 598048
rect 331218 597992 331274 598048
rect 331342 597992 331398 598048
rect 330970 597868 331026 597924
rect 331094 597868 331150 597924
rect 331218 597868 331274 597924
rect 331342 597868 331398 597924
rect 330970 597744 331026 597800
rect 331094 597744 331150 597800
rect 331218 597744 331274 597800
rect 331342 597744 331398 597800
rect 330970 586294 331026 586350
rect 331094 586294 331150 586350
rect 331218 586294 331274 586350
rect 331342 586294 331398 586350
rect 330970 586170 331026 586226
rect 331094 586170 331150 586226
rect 331218 586170 331274 586226
rect 331342 586170 331398 586226
rect 330970 586046 331026 586102
rect 331094 586046 331150 586102
rect 331218 586046 331274 586102
rect 331342 586046 331398 586102
rect 330970 585922 331026 585978
rect 331094 585922 331150 585978
rect 331218 585922 331274 585978
rect 331342 585922 331398 585978
rect 330970 568294 331026 568350
rect 331094 568294 331150 568350
rect 331218 568294 331274 568350
rect 331342 568294 331398 568350
rect 330970 568170 331026 568226
rect 331094 568170 331150 568226
rect 331218 568170 331274 568226
rect 331342 568170 331398 568226
rect 330970 568046 331026 568102
rect 331094 568046 331150 568102
rect 331218 568046 331274 568102
rect 331342 568046 331398 568102
rect 330970 567922 331026 567978
rect 331094 567922 331150 567978
rect 331218 567922 331274 567978
rect 331342 567922 331398 567978
rect 330970 550294 331026 550350
rect 331094 550294 331150 550350
rect 331218 550294 331274 550350
rect 331342 550294 331398 550350
rect 330970 550170 331026 550226
rect 331094 550170 331150 550226
rect 331218 550170 331274 550226
rect 331342 550170 331398 550226
rect 330970 550046 331026 550102
rect 331094 550046 331150 550102
rect 331218 550046 331274 550102
rect 331342 550046 331398 550102
rect 330970 549922 331026 549978
rect 331094 549922 331150 549978
rect 331218 549922 331274 549978
rect 331342 549922 331398 549978
rect 330970 532294 331026 532350
rect 331094 532294 331150 532350
rect 331218 532294 331274 532350
rect 331342 532294 331398 532350
rect 330970 532170 331026 532226
rect 331094 532170 331150 532226
rect 331218 532170 331274 532226
rect 331342 532170 331398 532226
rect 330970 532046 331026 532102
rect 331094 532046 331150 532102
rect 331218 532046 331274 532102
rect 331342 532046 331398 532102
rect 330970 531922 331026 531978
rect 331094 531922 331150 531978
rect 331218 531922 331274 531978
rect 331342 531922 331398 531978
rect 345250 597156 345306 597212
rect 345374 597156 345430 597212
rect 345498 597156 345554 597212
rect 345622 597156 345678 597212
rect 345250 597032 345306 597088
rect 345374 597032 345430 597088
rect 345498 597032 345554 597088
rect 345622 597032 345678 597088
rect 345250 596908 345306 596964
rect 345374 596908 345430 596964
rect 345498 596908 345554 596964
rect 345622 596908 345678 596964
rect 345250 596784 345306 596840
rect 345374 596784 345430 596840
rect 345498 596784 345554 596840
rect 345622 596784 345678 596840
rect 345250 580294 345306 580350
rect 345374 580294 345430 580350
rect 345498 580294 345554 580350
rect 345622 580294 345678 580350
rect 345250 580170 345306 580226
rect 345374 580170 345430 580226
rect 345498 580170 345554 580226
rect 345622 580170 345678 580226
rect 345250 580046 345306 580102
rect 345374 580046 345430 580102
rect 345498 580046 345554 580102
rect 345622 580046 345678 580102
rect 345250 579922 345306 579978
rect 345374 579922 345430 579978
rect 345498 579922 345554 579978
rect 345622 579922 345678 579978
rect 345250 562294 345306 562350
rect 345374 562294 345430 562350
rect 345498 562294 345554 562350
rect 345622 562294 345678 562350
rect 345250 562170 345306 562226
rect 345374 562170 345430 562226
rect 345498 562170 345554 562226
rect 345622 562170 345678 562226
rect 345250 562046 345306 562102
rect 345374 562046 345430 562102
rect 345498 562046 345554 562102
rect 345622 562046 345678 562102
rect 345250 561922 345306 561978
rect 345374 561922 345430 561978
rect 345498 561922 345554 561978
rect 345622 561922 345678 561978
rect 345250 544294 345306 544350
rect 345374 544294 345430 544350
rect 345498 544294 345554 544350
rect 345622 544294 345678 544350
rect 345250 544170 345306 544226
rect 345374 544170 345430 544226
rect 345498 544170 345554 544226
rect 345622 544170 345678 544226
rect 345250 544046 345306 544102
rect 345374 544046 345430 544102
rect 345498 544046 345554 544102
rect 345622 544046 345678 544102
rect 345250 543922 345306 543978
rect 345374 543922 345430 543978
rect 345498 543922 345554 543978
rect 345622 543922 345678 543978
rect 345250 526294 345306 526350
rect 345374 526294 345430 526350
rect 345498 526294 345554 526350
rect 345622 526294 345678 526350
rect 345250 526170 345306 526226
rect 345374 526170 345430 526226
rect 345498 526170 345554 526226
rect 345622 526170 345678 526226
rect 345250 526046 345306 526102
rect 345374 526046 345430 526102
rect 345498 526046 345554 526102
rect 345622 526046 345678 526102
rect 345250 525922 345306 525978
rect 345374 525922 345430 525978
rect 345498 525922 345554 525978
rect 345622 525922 345678 525978
rect 348970 598116 349026 598172
rect 349094 598116 349150 598172
rect 349218 598116 349274 598172
rect 349342 598116 349398 598172
rect 348970 597992 349026 598048
rect 349094 597992 349150 598048
rect 349218 597992 349274 598048
rect 349342 597992 349398 598048
rect 348970 597868 349026 597924
rect 349094 597868 349150 597924
rect 349218 597868 349274 597924
rect 349342 597868 349398 597924
rect 348970 597744 349026 597800
rect 349094 597744 349150 597800
rect 349218 597744 349274 597800
rect 349342 597744 349398 597800
rect 348970 586294 349026 586350
rect 349094 586294 349150 586350
rect 349218 586294 349274 586350
rect 349342 586294 349398 586350
rect 348970 586170 349026 586226
rect 349094 586170 349150 586226
rect 349218 586170 349274 586226
rect 349342 586170 349398 586226
rect 348970 586046 349026 586102
rect 349094 586046 349150 586102
rect 349218 586046 349274 586102
rect 349342 586046 349398 586102
rect 348970 585922 349026 585978
rect 349094 585922 349150 585978
rect 349218 585922 349274 585978
rect 349342 585922 349398 585978
rect 348970 568294 349026 568350
rect 349094 568294 349150 568350
rect 349218 568294 349274 568350
rect 349342 568294 349398 568350
rect 348970 568170 349026 568226
rect 349094 568170 349150 568226
rect 349218 568170 349274 568226
rect 349342 568170 349398 568226
rect 348970 568046 349026 568102
rect 349094 568046 349150 568102
rect 349218 568046 349274 568102
rect 349342 568046 349398 568102
rect 348970 567922 349026 567978
rect 349094 567922 349150 567978
rect 349218 567922 349274 567978
rect 349342 567922 349398 567978
rect 348970 550294 349026 550350
rect 349094 550294 349150 550350
rect 349218 550294 349274 550350
rect 349342 550294 349398 550350
rect 348970 550170 349026 550226
rect 349094 550170 349150 550226
rect 349218 550170 349274 550226
rect 349342 550170 349398 550226
rect 348970 550046 349026 550102
rect 349094 550046 349150 550102
rect 349218 550046 349274 550102
rect 349342 550046 349398 550102
rect 348970 549922 349026 549978
rect 349094 549922 349150 549978
rect 349218 549922 349274 549978
rect 349342 549922 349398 549978
rect 348970 532294 349026 532350
rect 349094 532294 349150 532350
rect 349218 532294 349274 532350
rect 349342 532294 349398 532350
rect 348970 532170 349026 532226
rect 349094 532170 349150 532226
rect 349218 532170 349274 532226
rect 349342 532170 349398 532226
rect 348970 532046 349026 532102
rect 349094 532046 349150 532102
rect 349218 532046 349274 532102
rect 349342 532046 349398 532102
rect 348970 531922 349026 531978
rect 349094 531922 349150 531978
rect 349218 531922 349274 531978
rect 349342 531922 349398 531978
rect 363250 597156 363306 597212
rect 363374 597156 363430 597212
rect 363498 597156 363554 597212
rect 363622 597156 363678 597212
rect 363250 597032 363306 597088
rect 363374 597032 363430 597088
rect 363498 597032 363554 597088
rect 363622 597032 363678 597088
rect 363250 596908 363306 596964
rect 363374 596908 363430 596964
rect 363498 596908 363554 596964
rect 363622 596908 363678 596964
rect 363250 596784 363306 596840
rect 363374 596784 363430 596840
rect 363498 596784 363554 596840
rect 363622 596784 363678 596840
rect 363250 580294 363306 580350
rect 363374 580294 363430 580350
rect 363498 580294 363554 580350
rect 363622 580294 363678 580350
rect 363250 580170 363306 580226
rect 363374 580170 363430 580226
rect 363498 580170 363554 580226
rect 363622 580170 363678 580226
rect 363250 580046 363306 580102
rect 363374 580046 363430 580102
rect 363498 580046 363554 580102
rect 363622 580046 363678 580102
rect 363250 579922 363306 579978
rect 363374 579922 363430 579978
rect 363498 579922 363554 579978
rect 363622 579922 363678 579978
rect 363250 562294 363306 562350
rect 363374 562294 363430 562350
rect 363498 562294 363554 562350
rect 363622 562294 363678 562350
rect 363250 562170 363306 562226
rect 363374 562170 363430 562226
rect 363498 562170 363554 562226
rect 363622 562170 363678 562226
rect 363250 562046 363306 562102
rect 363374 562046 363430 562102
rect 363498 562046 363554 562102
rect 363622 562046 363678 562102
rect 363250 561922 363306 561978
rect 363374 561922 363430 561978
rect 363498 561922 363554 561978
rect 363622 561922 363678 561978
rect 363250 544294 363306 544350
rect 363374 544294 363430 544350
rect 363498 544294 363554 544350
rect 363622 544294 363678 544350
rect 363250 544170 363306 544226
rect 363374 544170 363430 544226
rect 363498 544170 363554 544226
rect 363622 544170 363678 544226
rect 363250 544046 363306 544102
rect 363374 544046 363430 544102
rect 363498 544046 363554 544102
rect 363622 544046 363678 544102
rect 363250 543922 363306 543978
rect 363374 543922 363430 543978
rect 363498 543922 363554 543978
rect 363622 543922 363678 543978
rect 363250 526294 363306 526350
rect 363374 526294 363430 526350
rect 363498 526294 363554 526350
rect 363622 526294 363678 526350
rect 363250 526170 363306 526226
rect 363374 526170 363430 526226
rect 363498 526170 363554 526226
rect 363622 526170 363678 526226
rect 363250 526046 363306 526102
rect 363374 526046 363430 526102
rect 363498 526046 363554 526102
rect 363622 526046 363678 526102
rect 363250 525922 363306 525978
rect 363374 525922 363430 525978
rect 363498 525922 363554 525978
rect 363622 525922 363678 525978
rect 366970 598116 367026 598172
rect 367094 598116 367150 598172
rect 367218 598116 367274 598172
rect 367342 598116 367398 598172
rect 366970 597992 367026 598048
rect 367094 597992 367150 598048
rect 367218 597992 367274 598048
rect 367342 597992 367398 598048
rect 366970 597868 367026 597924
rect 367094 597868 367150 597924
rect 367218 597868 367274 597924
rect 367342 597868 367398 597924
rect 366970 597744 367026 597800
rect 367094 597744 367150 597800
rect 367218 597744 367274 597800
rect 367342 597744 367398 597800
rect 366970 586294 367026 586350
rect 367094 586294 367150 586350
rect 367218 586294 367274 586350
rect 367342 586294 367398 586350
rect 366970 586170 367026 586226
rect 367094 586170 367150 586226
rect 367218 586170 367274 586226
rect 367342 586170 367398 586226
rect 366970 586046 367026 586102
rect 367094 586046 367150 586102
rect 367218 586046 367274 586102
rect 367342 586046 367398 586102
rect 366970 585922 367026 585978
rect 367094 585922 367150 585978
rect 367218 585922 367274 585978
rect 367342 585922 367398 585978
rect 366970 568294 367026 568350
rect 367094 568294 367150 568350
rect 367218 568294 367274 568350
rect 367342 568294 367398 568350
rect 366970 568170 367026 568226
rect 367094 568170 367150 568226
rect 367218 568170 367274 568226
rect 367342 568170 367398 568226
rect 366970 568046 367026 568102
rect 367094 568046 367150 568102
rect 367218 568046 367274 568102
rect 367342 568046 367398 568102
rect 366970 567922 367026 567978
rect 367094 567922 367150 567978
rect 367218 567922 367274 567978
rect 367342 567922 367398 567978
rect 366970 550294 367026 550350
rect 367094 550294 367150 550350
rect 367218 550294 367274 550350
rect 367342 550294 367398 550350
rect 366970 550170 367026 550226
rect 367094 550170 367150 550226
rect 367218 550170 367274 550226
rect 367342 550170 367398 550226
rect 366970 550046 367026 550102
rect 367094 550046 367150 550102
rect 367218 550046 367274 550102
rect 367342 550046 367398 550102
rect 366970 549922 367026 549978
rect 367094 549922 367150 549978
rect 367218 549922 367274 549978
rect 367342 549922 367398 549978
rect 366970 532294 367026 532350
rect 367094 532294 367150 532350
rect 367218 532294 367274 532350
rect 367342 532294 367398 532350
rect 366970 532170 367026 532226
rect 367094 532170 367150 532226
rect 367218 532170 367274 532226
rect 367342 532170 367398 532226
rect 366970 532046 367026 532102
rect 367094 532046 367150 532102
rect 367218 532046 367274 532102
rect 367342 532046 367398 532102
rect 366970 531922 367026 531978
rect 367094 531922 367150 531978
rect 367218 531922 367274 531978
rect 367342 531922 367398 531978
rect 381250 597156 381306 597212
rect 381374 597156 381430 597212
rect 381498 597156 381554 597212
rect 381622 597156 381678 597212
rect 381250 597032 381306 597088
rect 381374 597032 381430 597088
rect 381498 597032 381554 597088
rect 381622 597032 381678 597088
rect 381250 596908 381306 596964
rect 381374 596908 381430 596964
rect 381498 596908 381554 596964
rect 381622 596908 381678 596964
rect 381250 596784 381306 596840
rect 381374 596784 381430 596840
rect 381498 596784 381554 596840
rect 381622 596784 381678 596840
rect 381250 580294 381306 580350
rect 381374 580294 381430 580350
rect 381498 580294 381554 580350
rect 381622 580294 381678 580350
rect 381250 580170 381306 580226
rect 381374 580170 381430 580226
rect 381498 580170 381554 580226
rect 381622 580170 381678 580226
rect 381250 580046 381306 580102
rect 381374 580046 381430 580102
rect 381498 580046 381554 580102
rect 381622 580046 381678 580102
rect 381250 579922 381306 579978
rect 381374 579922 381430 579978
rect 381498 579922 381554 579978
rect 381622 579922 381678 579978
rect 381250 562294 381306 562350
rect 381374 562294 381430 562350
rect 381498 562294 381554 562350
rect 381622 562294 381678 562350
rect 381250 562170 381306 562226
rect 381374 562170 381430 562226
rect 381498 562170 381554 562226
rect 381622 562170 381678 562226
rect 381250 562046 381306 562102
rect 381374 562046 381430 562102
rect 381498 562046 381554 562102
rect 381622 562046 381678 562102
rect 381250 561922 381306 561978
rect 381374 561922 381430 561978
rect 381498 561922 381554 561978
rect 381622 561922 381678 561978
rect 381250 544294 381306 544350
rect 381374 544294 381430 544350
rect 381498 544294 381554 544350
rect 381622 544294 381678 544350
rect 381250 544170 381306 544226
rect 381374 544170 381430 544226
rect 381498 544170 381554 544226
rect 381622 544170 381678 544226
rect 381250 544046 381306 544102
rect 381374 544046 381430 544102
rect 381498 544046 381554 544102
rect 381622 544046 381678 544102
rect 381250 543922 381306 543978
rect 381374 543922 381430 543978
rect 381498 543922 381554 543978
rect 381622 543922 381678 543978
rect 381250 526294 381306 526350
rect 381374 526294 381430 526350
rect 381498 526294 381554 526350
rect 381622 526294 381678 526350
rect 381250 526170 381306 526226
rect 381374 526170 381430 526226
rect 381498 526170 381554 526226
rect 381622 526170 381678 526226
rect 381250 526046 381306 526102
rect 381374 526046 381430 526102
rect 381498 526046 381554 526102
rect 381622 526046 381678 526102
rect 381250 525922 381306 525978
rect 381374 525922 381430 525978
rect 381498 525922 381554 525978
rect 381622 525922 381678 525978
rect 384970 598116 385026 598172
rect 385094 598116 385150 598172
rect 385218 598116 385274 598172
rect 385342 598116 385398 598172
rect 384970 597992 385026 598048
rect 385094 597992 385150 598048
rect 385218 597992 385274 598048
rect 385342 597992 385398 598048
rect 384970 597868 385026 597924
rect 385094 597868 385150 597924
rect 385218 597868 385274 597924
rect 385342 597868 385398 597924
rect 384970 597744 385026 597800
rect 385094 597744 385150 597800
rect 385218 597744 385274 597800
rect 385342 597744 385398 597800
rect 384970 586294 385026 586350
rect 385094 586294 385150 586350
rect 385218 586294 385274 586350
rect 385342 586294 385398 586350
rect 384970 586170 385026 586226
rect 385094 586170 385150 586226
rect 385218 586170 385274 586226
rect 385342 586170 385398 586226
rect 384970 586046 385026 586102
rect 385094 586046 385150 586102
rect 385218 586046 385274 586102
rect 385342 586046 385398 586102
rect 384970 585922 385026 585978
rect 385094 585922 385150 585978
rect 385218 585922 385274 585978
rect 385342 585922 385398 585978
rect 384970 568294 385026 568350
rect 385094 568294 385150 568350
rect 385218 568294 385274 568350
rect 385342 568294 385398 568350
rect 384970 568170 385026 568226
rect 385094 568170 385150 568226
rect 385218 568170 385274 568226
rect 385342 568170 385398 568226
rect 384970 568046 385026 568102
rect 385094 568046 385150 568102
rect 385218 568046 385274 568102
rect 385342 568046 385398 568102
rect 384970 567922 385026 567978
rect 385094 567922 385150 567978
rect 385218 567922 385274 567978
rect 385342 567922 385398 567978
rect 384970 550294 385026 550350
rect 385094 550294 385150 550350
rect 385218 550294 385274 550350
rect 385342 550294 385398 550350
rect 384970 550170 385026 550226
rect 385094 550170 385150 550226
rect 385218 550170 385274 550226
rect 385342 550170 385398 550226
rect 384970 550046 385026 550102
rect 385094 550046 385150 550102
rect 385218 550046 385274 550102
rect 385342 550046 385398 550102
rect 384970 549922 385026 549978
rect 385094 549922 385150 549978
rect 385218 549922 385274 549978
rect 385342 549922 385398 549978
rect 384970 532294 385026 532350
rect 385094 532294 385150 532350
rect 385218 532294 385274 532350
rect 385342 532294 385398 532350
rect 384970 532170 385026 532226
rect 385094 532170 385150 532226
rect 385218 532170 385274 532226
rect 385342 532170 385398 532226
rect 384970 532046 385026 532102
rect 385094 532046 385150 532102
rect 385218 532046 385274 532102
rect 385342 532046 385398 532102
rect 384970 531922 385026 531978
rect 385094 531922 385150 531978
rect 385218 531922 385274 531978
rect 385342 531922 385398 531978
rect 399250 597156 399306 597212
rect 399374 597156 399430 597212
rect 399498 597156 399554 597212
rect 399622 597156 399678 597212
rect 399250 597032 399306 597088
rect 399374 597032 399430 597088
rect 399498 597032 399554 597088
rect 399622 597032 399678 597088
rect 399250 596908 399306 596964
rect 399374 596908 399430 596964
rect 399498 596908 399554 596964
rect 399622 596908 399678 596964
rect 399250 596784 399306 596840
rect 399374 596784 399430 596840
rect 399498 596784 399554 596840
rect 399622 596784 399678 596840
rect 399250 580294 399306 580350
rect 399374 580294 399430 580350
rect 399498 580294 399554 580350
rect 399622 580294 399678 580350
rect 399250 580170 399306 580226
rect 399374 580170 399430 580226
rect 399498 580170 399554 580226
rect 399622 580170 399678 580226
rect 399250 580046 399306 580102
rect 399374 580046 399430 580102
rect 399498 580046 399554 580102
rect 399622 580046 399678 580102
rect 399250 579922 399306 579978
rect 399374 579922 399430 579978
rect 399498 579922 399554 579978
rect 399622 579922 399678 579978
rect 399250 562294 399306 562350
rect 399374 562294 399430 562350
rect 399498 562294 399554 562350
rect 399622 562294 399678 562350
rect 399250 562170 399306 562226
rect 399374 562170 399430 562226
rect 399498 562170 399554 562226
rect 399622 562170 399678 562226
rect 399250 562046 399306 562102
rect 399374 562046 399430 562102
rect 399498 562046 399554 562102
rect 399622 562046 399678 562102
rect 399250 561922 399306 561978
rect 399374 561922 399430 561978
rect 399498 561922 399554 561978
rect 399622 561922 399678 561978
rect 399250 544294 399306 544350
rect 399374 544294 399430 544350
rect 399498 544294 399554 544350
rect 399622 544294 399678 544350
rect 399250 544170 399306 544226
rect 399374 544170 399430 544226
rect 399498 544170 399554 544226
rect 399622 544170 399678 544226
rect 399250 544046 399306 544102
rect 399374 544046 399430 544102
rect 399498 544046 399554 544102
rect 399622 544046 399678 544102
rect 399250 543922 399306 543978
rect 399374 543922 399430 543978
rect 399498 543922 399554 543978
rect 399622 543922 399678 543978
rect 399250 526294 399306 526350
rect 399374 526294 399430 526350
rect 399498 526294 399554 526350
rect 399622 526294 399678 526350
rect 399250 526170 399306 526226
rect 399374 526170 399430 526226
rect 399498 526170 399554 526226
rect 399622 526170 399678 526226
rect 399250 526046 399306 526102
rect 399374 526046 399430 526102
rect 399498 526046 399554 526102
rect 399622 526046 399678 526102
rect 399250 525922 399306 525978
rect 399374 525922 399430 525978
rect 399498 525922 399554 525978
rect 399622 525922 399678 525978
rect 402970 598116 403026 598172
rect 403094 598116 403150 598172
rect 403218 598116 403274 598172
rect 403342 598116 403398 598172
rect 402970 597992 403026 598048
rect 403094 597992 403150 598048
rect 403218 597992 403274 598048
rect 403342 597992 403398 598048
rect 402970 597868 403026 597924
rect 403094 597868 403150 597924
rect 403218 597868 403274 597924
rect 403342 597868 403398 597924
rect 402970 597744 403026 597800
rect 403094 597744 403150 597800
rect 403218 597744 403274 597800
rect 403342 597744 403398 597800
rect 402970 586294 403026 586350
rect 403094 586294 403150 586350
rect 403218 586294 403274 586350
rect 403342 586294 403398 586350
rect 402970 586170 403026 586226
rect 403094 586170 403150 586226
rect 403218 586170 403274 586226
rect 403342 586170 403398 586226
rect 402970 586046 403026 586102
rect 403094 586046 403150 586102
rect 403218 586046 403274 586102
rect 403342 586046 403398 586102
rect 402970 585922 403026 585978
rect 403094 585922 403150 585978
rect 403218 585922 403274 585978
rect 403342 585922 403398 585978
rect 402970 568294 403026 568350
rect 403094 568294 403150 568350
rect 403218 568294 403274 568350
rect 403342 568294 403398 568350
rect 402970 568170 403026 568226
rect 403094 568170 403150 568226
rect 403218 568170 403274 568226
rect 403342 568170 403398 568226
rect 402970 568046 403026 568102
rect 403094 568046 403150 568102
rect 403218 568046 403274 568102
rect 403342 568046 403398 568102
rect 402970 567922 403026 567978
rect 403094 567922 403150 567978
rect 403218 567922 403274 567978
rect 403342 567922 403398 567978
rect 402970 550294 403026 550350
rect 403094 550294 403150 550350
rect 403218 550294 403274 550350
rect 403342 550294 403398 550350
rect 402970 550170 403026 550226
rect 403094 550170 403150 550226
rect 403218 550170 403274 550226
rect 403342 550170 403398 550226
rect 402970 550046 403026 550102
rect 403094 550046 403150 550102
rect 403218 550046 403274 550102
rect 403342 550046 403398 550102
rect 402970 549922 403026 549978
rect 403094 549922 403150 549978
rect 403218 549922 403274 549978
rect 403342 549922 403398 549978
rect 402970 532294 403026 532350
rect 403094 532294 403150 532350
rect 403218 532294 403274 532350
rect 403342 532294 403398 532350
rect 402970 532170 403026 532226
rect 403094 532170 403150 532226
rect 403218 532170 403274 532226
rect 403342 532170 403398 532226
rect 402970 532046 403026 532102
rect 403094 532046 403150 532102
rect 403218 532046 403274 532102
rect 403342 532046 403398 532102
rect 402970 531922 403026 531978
rect 403094 531922 403150 531978
rect 403218 531922 403274 531978
rect 403342 531922 403398 531978
rect 417250 597156 417306 597212
rect 417374 597156 417430 597212
rect 417498 597156 417554 597212
rect 417622 597156 417678 597212
rect 417250 597032 417306 597088
rect 417374 597032 417430 597088
rect 417498 597032 417554 597088
rect 417622 597032 417678 597088
rect 417250 596908 417306 596964
rect 417374 596908 417430 596964
rect 417498 596908 417554 596964
rect 417622 596908 417678 596964
rect 417250 596784 417306 596840
rect 417374 596784 417430 596840
rect 417498 596784 417554 596840
rect 417622 596784 417678 596840
rect 417250 580294 417306 580350
rect 417374 580294 417430 580350
rect 417498 580294 417554 580350
rect 417622 580294 417678 580350
rect 417250 580170 417306 580226
rect 417374 580170 417430 580226
rect 417498 580170 417554 580226
rect 417622 580170 417678 580226
rect 417250 580046 417306 580102
rect 417374 580046 417430 580102
rect 417498 580046 417554 580102
rect 417622 580046 417678 580102
rect 417250 579922 417306 579978
rect 417374 579922 417430 579978
rect 417498 579922 417554 579978
rect 417622 579922 417678 579978
rect 417250 562294 417306 562350
rect 417374 562294 417430 562350
rect 417498 562294 417554 562350
rect 417622 562294 417678 562350
rect 417250 562170 417306 562226
rect 417374 562170 417430 562226
rect 417498 562170 417554 562226
rect 417622 562170 417678 562226
rect 417250 562046 417306 562102
rect 417374 562046 417430 562102
rect 417498 562046 417554 562102
rect 417622 562046 417678 562102
rect 417250 561922 417306 561978
rect 417374 561922 417430 561978
rect 417498 561922 417554 561978
rect 417622 561922 417678 561978
rect 417250 544294 417306 544350
rect 417374 544294 417430 544350
rect 417498 544294 417554 544350
rect 417622 544294 417678 544350
rect 417250 544170 417306 544226
rect 417374 544170 417430 544226
rect 417498 544170 417554 544226
rect 417622 544170 417678 544226
rect 417250 544046 417306 544102
rect 417374 544046 417430 544102
rect 417498 544046 417554 544102
rect 417622 544046 417678 544102
rect 417250 543922 417306 543978
rect 417374 543922 417430 543978
rect 417498 543922 417554 543978
rect 417622 543922 417678 543978
rect 417250 526294 417306 526350
rect 417374 526294 417430 526350
rect 417498 526294 417554 526350
rect 417622 526294 417678 526350
rect 417250 526170 417306 526226
rect 417374 526170 417430 526226
rect 417498 526170 417554 526226
rect 417622 526170 417678 526226
rect 417250 526046 417306 526102
rect 417374 526046 417430 526102
rect 417498 526046 417554 526102
rect 417622 526046 417678 526102
rect 417250 525922 417306 525978
rect 417374 525922 417430 525978
rect 417498 525922 417554 525978
rect 417622 525922 417678 525978
rect 420970 598116 421026 598172
rect 421094 598116 421150 598172
rect 421218 598116 421274 598172
rect 421342 598116 421398 598172
rect 420970 597992 421026 598048
rect 421094 597992 421150 598048
rect 421218 597992 421274 598048
rect 421342 597992 421398 598048
rect 420970 597868 421026 597924
rect 421094 597868 421150 597924
rect 421218 597868 421274 597924
rect 421342 597868 421398 597924
rect 420970 597744 421026 597800
rect 421094 597744 421150 597800
rect 421218 597744 421274 597800
rect 421342 597744 421398 597800
rect 420970 586294 421026 586350
rect 421094 586294 421150 586350
rect 421218 586294 421274 586350
rect 421342 586294 421398 586350
rect 420970 586170 421026 586226
rect 421094 586170 421150 586226
rect 421218 586170 421274 586226
rect 421342 586170 421398 586226
rect 420970 586046 421026 586102
rect 421094 586046 421150 586102
rect 421218 586046 421274 586102
rect 421342 586046 421398 586102
rect 420970 585922 421026 585978
rect 421094 585922 421150 585978
rect 421218 585922 421274 585978
rect 421342 585922 421398 585978
rect 420970 568294 421026 568350
rect 421094 568294 421150 568350
rect 421218 568294 421274 568350
rect 421342 568294 421398 568350
rect 420970 568170 421026 568226
rect 421094 568170 421150 568226
rect 421218 568170 421274 568226
rect 421342 568170 421398 568226
rect 420970 568046 421026 568102
rect 421094 568046 421150 568102
rect 421218 568046 421274 568102
rect 421342 568046 421398 568102
rect 420970 567922 421026 567978
rect 421094 567922 421150 567978
rect 421218 567922 421274 567978
rect 421342 567922 421398 567978
rect 420970 550294 421026 550350
rect 421094 550294 421150 550350
rect 421218 550294 421274 550350
rect 421342 550294 421398 550350
rect 420970 550170 421026 550226
rect 421094 550170 421150 550226
rect 421218 550170 421274 550226
rect 421342 550170 421398 550226
rect 420970 550046 421026 550102
rect 421094 550046 421150 550102
rect 421218 550046 421274 550102
rect 421342 550046 421398 550102
rect 420970 549922 421026 549978
rect 421094 549922 421150 549978
rect 421218 549922 421274 549978
rect 421342 549922 421398 549978
rect 420970 532294 421026 532350
rect 421094 532294 421150 532350
rect 421218 532294 421274 532350
rect 421342 532294 421398 532350
rect 420970 532170 421026 532226
rect 421094 532170 421150 532226
rect 421218 532170 421274 532226
rect 421342 532170 421398 532226
rect 420970 532046 421026 532102
rect 421094 532046 421150 532102
rect 421218 532046 421274 532102
rect 421342 532046 421398 532102
rect 420970 531922 421026 531978
rect 421094 531922 421150 531978
rect 421218 531922 421274 531978
rect 421342 531922 421398 531978
rect 435250 597156 435306 597212
rect 435374 597156 435430 597212
rect 435498 597156 435554 597212
rect 435622 597156 435678 597212
rect 435250 597032 435306 597088
rect 435374 597032 435430 597088
rect 435498 597032 435554 597088
rect 435622 597032 435678 597088
rect 435250 596908 435306 596964
rect 435374 596908 435430 596964
rect 435498 596908 435554 596964
rect 435622 596908 435678 596964
rect 435250 596784 435306 596840
rect 435374 596784 435430 596840
rect 435498 596784 435554 596840
rect 435622 596784 435678 596840
rect 435250 580294 435306 580350
rect 435374 580294 435430 580350
rect 435498 580294 435554 580350
rect 435622 580294 435678 580350
rect 435250 580170 435306 580226
rect 435374 580170 435430 580226
rect 435498 580170 435554 580226
rect 435622 580170 435678 580226
rect 435250 580046 435306 580102
rect 435374 580046 435430 580102
rect 435498 580046 435554 580102
rect 435622 580046 435678 580102
rect 435250 579922 435306 579978
rect 435374 579922 435430 579978
rect 435498 579922 435554 579978
rect 435622 579922 435678 579978
rect 435250 562294 435306 562350
rect 435374 562294 435430 562350
rect 435498 562294 435554 562350
rect 435622 562294 435678 562350
rect 435250 562170 435306 562226
rect 435374 562170 435430 562226
rect 435498 562170 435554 562226
rect 435622 562170 435678 562226
rect 435250 562046 435306 562102
rect 435374 562046 435430 562102
rect 435498 562046 435554 562102
rect 435622 562046 435678 562102
rect 435250 561922 435306 561978
rect 435374 561922 435430 561978
rect 435498 561922 435554 561978
rect 435622 561922 435678 561978
rect 435250 544294 435306 544350
rect 435374 544294 435430 544350
rect 435498 544294 435554 544350
rect 435622 544294 435678 544350
rect 435250 544170 435306 544226
rect 435374 544170 435430 544226
rect 435498 544170 435554 544226
rect 435622 544170 435678 544226
rect 435250 544046 435306 544102
rect 435374 544046 435430 544102
rect 435498 544046 435554 544102
rect 435622 544046 435678 544102
rect 435250 543922 435306 543978
rect 435374 543922 435430 543978
rect 435498 543922 435554 543978
rect 435622 543922 435678 543978
rect 435250 526294 435306 526350
rect 435374 526294 435430 526350
rect 435498 526294 435554 526350
rect 435622 526294 435678 526350
rect 435250 526170 435306 526226
rect 435374 526170 435430 526226
rect 435498 526170 435554 526226
rect 435622 526170 435678 526226
rect 435250 526046 435306 526102
rect 435374 526046 435430 526102
rect 435498 526046 435554 526102
rect 435622 526046 435678 526102
rect 435250 525922 435306 525978
rect 435374 525922 435430 525978
rect 435498 525922 435554 525978
rect 435622 525922 435678 525978
rect 438970 598116 439026 598172
rect 439094 598116 439150 598172
rect 439218 598116 439274 598172
rect 439342 598116 439398 598172
rect 438970 597992 439026 598048
rect 439094 597992 439150 598048
rect 439218 597992 439274 598048
rect 439342 597992 439398 598048
rect 438970 597868 439026 597924
rect 439094 597868 439150 597924
rect 439218 597868 439274 597924
rect 439342 597868 439398 597924
rect 438970 597744 439026 597800
rect 439094 597744 439150 597800
rect 439218 597744 439274 597800
rect 439342 597744 439398 597800
rect 438970 586294 439026 586350
rect 439094 586294 439150 586350
rect 439218 586294 439274 586350
rect 439342 586294 439398 586350
rect 438970 586170 439026 586226
rect 439094 586170 439150 586226
rect 439218 586170 439274 586226
rect 439342 586170 439398 586226
rect 438970 586046 439026 586102
rect 439094 586046 439150 586102
rect 439218 586046 439274 586102
rect 439342 586046 439398 586102
rect 438970 585922 439026 585978
rect 439094 585922 439150 585978
rect 439218 585922 439274 585978
rect 439342 585922 439398 585978
rect 438970 568294 439026 568350
rect 439094 568294 439150 568350
rect 439218 568294 439274 568350
rect 439342 568294 439398 568350
rect 438970 568170 439026 568226
rect 439094 568170 439150 568226
rect 439218 568170 439274 568226
rect 439342 568170 439398 568226
rect 438970 568046 439026 568102
rect 439094 568046 439150 568102
rect 439218 568046 439274 568102
rect 439342 568046 439398 568102
rect 438970 567922 439026 567978
rect 439094 567922 439150 567978
rect 439218 567922 439274 567978
rect 439342 567922 439398 567978
rect 438970 550294 439026 550350
rect 439094 550294 439150 550350
rect 439218 550294 439274 550350
rect 439342 550294 439398 550350
rect 438970 550170 439026 550226
rect 439094 550170 439150 550226
rect 439218 550170 439274 550226
rect 439342 550170 439398 550226
rect 438970 550046 439026 550102
rect 439094 550046 439150 550102
rect 439218 550046 439274 550102
rect 439342 550046 439398 550102
rect 438970 549922 439026 549978
rect 439094 549922 439150 549978
rect 439218 549922 439274 549978
rect 439342 549922 439398 549978
rect 438970 532294 439026 532350
rect 439094 532294 439150 532350
rect 439218 532294 439274 532350
rect 439342 532294 439398 532350
rect 438970 532170 439026 532226
rect 439094 532170 439150 532226
rect 439218 532170 439274 532226
rect 439342 532170 439398 532226
rect 438970 532046 439026 532102
rect 439094 532046 439150 532102
rect 439218 532046 439274 532102
rect 439342 532046 439398 532102
rect 438970 531922 439026 531978
rect 439094 531922 439150 531978
rect 439218 531922 439274 531978
rect 439342 531922 439398 531978
rect 453250 597156 453306 597212
rect 453374 597156 453430 597212
rect 453498 597156 453554 597212
rect 453622 597156 453678 597212
rect 453250 597032 453306 597088
rect 453374 597032 453430 597088
rect 453498 597032 453554 597088
rect 453622 597032 453678 597088
rect 453250 596908 453306 596964
rect 453374 596908 453430 596964
rect 453498 596908 453554 596964
rect 453622 596908 453678 596964
rect 453250 596784 453306 596840
rect 453374 596784 453430 596840
rect 453498 596784 453554 596840
rect 453622 596784 453678 596840
rect 453250 580294 453306 580350
rect 453374 580294 453430 580350
rect 453498 580294 453554 580350
rect 453622 580294 453678 580350
rect 453250 580170 453306 580226
rect 453374 580170 453430 580226
rect 453498 580170 453554 580226
rect 453622 580170 453678 580226
rect 453250 580046 453306 580102
rect 453374 580046 453430 580102
rect 453498 580046 453554 580102
rect 453622 580046 453678 580102
rect 453250 579922 453306 579978
rect 453374 579922 453430 579978
rect 453498 579922 453554 579978
rect 453622 579922 453678 579978
rect 453250 562294 453306 562350
rect 453374 562294 453430 562350
rect 453498 562294 453554 562350
rect 453622 562294 453678 562350
rect 453250 562170 453306 562226
rect 453374 562170 453430 562226
rect 453498 562170 453554 562226
rect 453622 562170 453678 562226
rect 453250 562046 453306 562102
rect 453374 562046 453430 562102
rect 453498 562046 453554 562102
rect 453622 562046 453678 562102
rect 453250 561922 453306 561978
rect 453374 561922 453430 561978
rect 453498 561922 453554 561978
rect 453622 561922 453678 561978
rect 453250 544294 453306 544350
rect 453374 544294 453430 544350
rect 453498 544294 453554 544350
rect 453622 544294 453678 544350
rect 453250 544170 453306 544226
rect 453374 544170 453430 544226
rect 453498 544170 453554 544226
rect 453622 544170 453678 544226
rect 453250 544046 453306 544102
rect 453374 544046 453430 544102
rect 453498 544046 453554 544102
rect 453622 544046 453678 544102
rect 453250 543922 453306 543978
rect 453374 543922 453430 543978
rect 453498 543922 453554 543978
rect 453622 543922 453678 543978
rect 453250 526294 453306 526350
rect 453374 526294 453430 526350
rect 453498 526294 453554 526350
rect 453622 526294 453678 526350
rect 453250 526170 453306 526226
rect 453374 526170 453430 526226
rect 453498 526170 453554 526226
rect 453622 526170 453678 526226
rect 453250 526046 453306 526102
rect 453374 526046 453430 526102
rect 453498 526046 453554 526102
rect 453622 526046 453678 526102
rect 453250 525922 453306 525978
rect 453374 525922 453430 525978
rect 453498 525922 453554 525978
rect 453622 525922 453678 525978
rect 456970 598116 457026 598172
rect 457094 598116 457150 598172
rect 457218 598116 457274 598172
rect 457342 598116 457398 598172
rect 456970 597992 457026 598048
rect 457094 597992 457150 598048
rect 457218 597992 457274 598048
rect 457342 597992 457398 598048
rect 456970 597868 457026 597924
rect 457094 597868 457150 597924
rect 457218 597868 457274 597924
rect 457342 597868 457398 597924
rect 456970 597744 457026 597800
rect 457094 597744 457150 597800
rect 457218 597744 457274 597800
rect 457342 597744 457398 597800
rect 456970 586294 457026 586350
rect 457094 586294 457150 586350
rect 457218 586294 457274 586350
rect 457342 586294 457398 586350
rect 456970 586170 457026 586226
rect 457094 586170 457150 586226
rect 457218 586170 457274 586226
rect 457342 586170 457398 586226
rect 456970 586046 457026 586102
rect 457094 586046 457150 586102
rect 457218 586046 457274 586102
rect 457342 586046 457398 586102
rect 456970 585922 457026 585978
rect 457094 585922 457150 585978
rect 457218 585922 457274 585978
rect 457342 585922 457398 585978
rect 456970 568294 457026 568350
rect 457094 568294 457150 568350
rect 457218 568294 457274 568350
rect 457342 568294 457398 568350
rect 456970 568170 457026 568226
rect 457094 568170 457150 568226
rect 457218 568170 457274 568226
rect 457342 568170 457398 568226
rect 456970 568046 457026 568102
rect 457094 568046 457150 568102
rect 457218 568046 457274 568102
rect 457342 568046 457398 568102
rect 456970 567922 457026 567978
rect 457094 567922 457150 567978
rect 457218 567922 457274 567978
rect 457342 567922 457398 567978
rect 456970 550294 457026 550350
rect 457094 550294 457150 550350
rect 457218 550294 457274 550350
rect 457342 550294 457398 550350
rect 456970 550170 457026 550226
rect 457094 550170 457150 550226
rect 457218 550170 457274 550226
rect 457342 550170 457398 550226
rect 456970 550046 457026 550102
rect 457094 550046 457150 550102
rect 457218 550046 457274 550102
rect 457342 550046 457398 550102
rect 456970 549922 457026 549978
rect 457094 549922 457150 549978
rect 457218 549922 457274 549978
rect 457342 549922 457398 549978
rect 456970 532294 457026 532350
rect 457094 532294 457150 532350
rect 457218 532294 457274 532350
rect 457342 532294 457398 532350
rect 456970 532170 457026 532226
rect 457094 532170 457150 532226
rect 457218 532170 457274 532226
rect 457342 532170 457398 532226
rect 456970 532046 457026 532102
rect 457094 532046 457150 532102
rect 457218 532046 457274 532102
rect 457342 532046 457398 532102
rect 456970 531922 457026 531978
rect 457094 531922 457150 531978
rect 457218 531922 457274 531978
rect 457342 531922 457398 531978
rect 471250 597156 471306 597212
rect 471374 597156 471430 597212
rect 471498 597156 471554 597212
rect 471622 597156 471678 597212
rect 471250 597032 471306 597088
rect 471374 597032 471430 597088
rect 471498 597032 471554 597088
rect 471622 597032 471678 597088
rect 471250 596908 471306 596964
rect 471374 596908 471430 596964
rect 471498 596908 471554 596964
rect 471622 596908 471678 596964
rect 471250 596784 471306 596840
rect 471374 596784 471430 596840
rect 471498 596784 471554 596840
rect 471622 596784 471678 596840
rect 471250 580294 471306 580350
rect 471374 580294 471430 580350
rect 471498 580294 471554 580350
rect 471622 580294 471678 580350
rect 471250 580170 471306 580226
rect 471374 580170 471430 580226
rect 471498 580170 471554 580226
rect 471622 580170 471678 580226
rect 471250 580046 471306 580102
rect 471374 580046 471430 580102
rect 471498 580046 471554 580102
rect 471622 580046 471678 580102
rect 471250 579922 471306 579978
rect 471374 579922 471430 579978
rect 471498 579922 471554 579978
rect 471622 579922 471678 579978
rect 471250 562294 471306 562350
rect 471374 562294 471430 562350
rect 471498 562294 471554 562350
rect 471622 562294 471678 562350
rect 471250 562170 471306 562226
rect 471374 562170 471430 562226
rect 471498 562170 471554 562226
rect 471622 562170 471678 562226
rect 471250 562046 471306 562102
rect 471374 562046 471430 562102
rect 471498 562046 471554 562102
rect 471622 562046 471678 562102
rect 471250 561922 471306 561978
rect 471374 561922 471430 561978
rect 471498 561922 471554 561978
rect 471622 561922 471678 561978
rect 471250 544294 471306 544350
rect 471374 544294 471430 544350
rect 471498 544294 471554 544350
rect 471622 544294 471678 544350
rect 471250 544170 471306 544226
rect 471374 544170 471430 544226
rect 471498 544170 471554 544226
rect 471622 544170 471678 544226
rect 471250 544046 471306 544102
rect 471374 544046 471430 544102
rect 471498 544046 471554 544102
rect 471622 544046 471678 544102
rect 471250 543922 471306 543978
rect 471374 543922 471430 543978
rect 471498 543922 471554 543978
rect 471622 543922 471678 543978
rect 471250 526294 471306 526350
rect 471374 526294 471430 526350
rect 471498 526294 471554 526350
rect 471622 526294 471678 526350
rect 471250 526170 471306 526226
rect 471374 526170 471430 526226
rect 471498 526170 471554 526226
rect 471622 526170 471678 526226
rect 471250 526046 471306 526102
rect 471374 526046 471430 526102
rect 471498 526046 471554 526102
rect 471622 526046 471678 526102
rect 471250 525922 471306 525978
rect 471374 525922 471430 525978
rect 471498 525922 471554 525978
rect 471622 525922 471678 525978
rect 474970 598116 475026 598172
rect 475094 598116 475150 598172
rect 475218 598116 475274 598172
rect 475342 598116 475398 598172
rect 474970 597992 475026 598048
rect 475094 597992 475150 598048
rect 475218 597992 475274 598048
rect 475342 597992 475398 598048
rect 474970 597868 475026 597924
rect 475094 597868 475150 597924
rect 475218 597868 475274 597924
rect 475342 597868 475398 597924
rect 474970 597744 475026 597800
rect 475094 597744 475150 597800
rect 475218 597744 475274 597800
rect 475342 597744 475398 597800
rect 474970 586294 475026 586350
rect 475094 586294 475150 586350
rect 475218 586294 475274 586350
rect 475342 586294 475398 586350
rect 474970 586170 475026 586226
rect 475094 586170 475150 586226
rect 475218 586170 475274 586226
rect 475342 586170 475398 586226
rect 474970 586046 475026 586102
rect 475094 586046 475150 586102
rect 475218 586046 475274 586102
rect 475342 586046 475398 586102
rect 474970 585922 475026 585978
rect 475094 585922 475150 585978
rect 475218 585922 475274 585978
rect 475342 585922 475398 585978
rect 474970 568294 475026 568350
rect 475094 568294 475150 568350
rect 475218 568294 475274 568350
rect 475342 568294 475398 568350
rect 474970 568170 475026 568226
rect 475094 568170 475150 568226
rect 475218 568170 475274 568226
rect 475342 568170 475398 568226
rect 474970 568046 475026 568102
rect 475094 568046 475150 568102
rect 475218 568046 475274 568102
rect 475342 568046 475398 568102
rect 474970 567922 475026 567978
rect 475094 567922 475150 567978
rect 475218 567922 475274 567978
rect 475342 567922 475398 567978
rect 474970 550294 475026 550350
rect 475094 550294 475150 550350
rect 475218 550294 475274 550350
rect 475342 550294 475398 550350
rect 474970 550170 475026 550226
rect 475094 550170 475150 550226
rect 475218 550170 475274 550226
rect 475342 550170 475398 550226
rect 474970 550046 475026 550102
rect 475094 550046 475150 550102
rect 475218 550046 475274 550102
rect 475342 550046 475398 550102
rect 474970 549922 475026 549978
rect 475094 549922 475150 549978
rect 475218 549922 475274 549978
rect 475342 549922 475398 549978
rect 474970 532294 475026 532350
rect 475094 532294 475150 532350
rect 475218 532294 475274 532350
rect 475342 532294 475398 532350
rect 474970 532170 475026 532226
rect 475094 532170 475150 532226
rect 475218 532170 475274 532226
rect 475342 532170 475398 532226
rect 474970 532046 475026 532102
rect 475094 532046 475150 532102
rect 475218 532046 475274 532102
rect 475342 532046 475398 532102
rect 474970 531922 475026 531978
rect 475094 531922 475150 531978
rect 475218 531922 475274 531978
rect 475342 531922 475398 531978
rect 489250 597156 489306 597212
rect 489374 597156 489430 597212
rect 489498 597156 489554 597212
rect 489622 597156 489678 597212
rect 489250 597032 489306 597088
rect 489374 597032 489430 597088
rect 489498 597032 489554 597088
rect 489622 597032 489678 597088
rect 489250 596908 489306 596964
rect 489374 596908 489430 596964
rect 489498 596908 489554 596964
rect 489622 596908 489678 596964
rect 489250 596784 489306 596840
rect 489374 596784 489430 596840
rect 489498 596784 489554 596840
rect 489622 596784 489678 596840
rect 489250 580294 489306 580350
rect 489374 580294 489430 580350
rect 489498 580294 489554 580350
rect 489622 580294 489678 580350
rect 489250 580170 489306 580226
rect 489374 580170 489430 580226
rect 489498 580170 489554 580226
rect 489622 580170 489678 580226
rect 489250 580046 489306 580102
rect 489374 580046 489430 580102
rect 489498 580046 489554 580102
rect 489622 580046 489678 580102
rect 489250 579922 489306 579978
rect 489374 579922 489430 579978
rect 489498 579922 489554 579978
rect 489622 579922 489678 579978
rect 489250 562294 489306 562350
rect 489374 562294 489430 562350
rect 489498 562294 489554 562350
rect 489622 562294 489678 562350
rect 489250 562170 489306 562226
rect 489374 562170 489430 562226
rect 489498 562170 489554 562226
rect 489622 562170 489678 562226
rect 489250 562046 489306 562102
rect 489374 562046 489430 562102
rect 489498 562046 489554 562102
rect 489622 562046 489678 562102
rect 489250 561922 489306 561978
rect 489374 561922 489430 561978
rect 489498 561922 489554 561978
rect 489622 561922 489678 561978
rect 489250 544294 489306 544350
rect 489374 544294 489430 544350
rect 489498 544294 489554 544350
rect 489622 544294 489678 544350
rect 489250 544170 489306 544226
rect 489374 544170 489430 544226
rect 489498 544170 489554 544226
rect 489622 544170 489678 544226
rect 489250 544046 489306 544102
rect 489374 544046 489430 544102
rect 489498 544046 489554 544102
rect 489622 544046 489678 544102
rect 489250 543922 489306 543978
rect 489374 543922 489430 543978
rect 489498 543922 489554 543978
rect 489622 543922 489678 543978
rect 489250 526294 489306 526350
rect 489374 526294 489430 526350
rect 489498 526294 489554 526350
rect 489622 526294 489678 526350
rect 489250 526170 489306 526226
rect 489374 526170 489430 526226
rect 489498 526170 489554 526226
rect 489622 526170 489678 526226
rect 489250 526046 489306 526102
rect 489374 526046 489430 526102
rect 489498 526046 489554 526102
rect 489622 526046 489678 526102
rect 489250 525922 489306 525978
rect 489374 525922 489430 525978
rect 489498 525922 489554 525978
rect 489622 525922 489678 525978
rect 492970 598116 493026 598172
rect 493094 598116 493150 598172
rect 493218 598116 493274 598172
rect 493342 598116 493398 598172
rect 492970 597992 493026 598048
rect 493094 597992 493150 598048
rect 493218 597992 493274 598048
rect 493342 597992 493398 598048
rect 492970 597868 493026 597924
rect 493094 597868 493150 597924
rect 493218 597868 493274 597924
rect 493342 597868 493398 597924
rect 492970 597744 493026 597800
rect 493094 597744 493150 597800
rect 493218 597744 493274 597800
rect 493342 597744 493398 597800
rect 492970 586294 493026 586350
rect 493094 586294 493150 586350
rect 493218 586294 493274 586350
rect 493342 586294 493398 586350
rect 492970 586170 493026 586226
rect 493094 586170 493150 586226
rect 493218 586170 493274 586226
rect 493342 586170 493398 586226
rect 492970 586046 493026 586102
rect 493094 586046 493150 586102
rect 493218 586046 493274 586102
rect 493342 586046 493398 586102
rect 492970 585922 493026 585978
rect 493094 585922 493150 585978
rect 493218 585922 493274 585978
rect 493342 585922 493398 585978
rect 492970 568294 493026 568350
rect 493094 568294 493150 568350
rect 493218 568294 493274 568350
rect 493342 568294 493398 568350
rect 492970 568170 493026 568226
rect 493094 568170 493150 568226
rect 493218 568170 493274 568226
rect 493342 568170 493398 568226
rect 492970 568046 493026 568102
rect 493094 568046 493150 568102
rect 493218 568046 493274 568102
rect 493342 568046 493398 568102
rect 492970 567922 493026 567978
rect 493094 567922 493150 567978
rect 493218 567922 493274 567978
rect 493342 567922 493398 567978
rect 492970 550294 493026 550350
rect 493094 550294 493150 550350
rect 493218 550294 493274 550350
rect 493342 550294 493398 550350
rect 492970 550170 493026 550226
rect 493094 550170 493150 550226
rect 493218 550170 493274 550226
rect 493342 550170 493398 550226
rect 492970 550046 493026 550102
rect 493094 550046 493150 550102
rect 493218 550046 493274 550102
rect 493342 550046 493398 550102
rect 492970 549922 493026 549978
rect 493094 549922 493150 549978
rect 493218 549922 493274 549978
rect 493342 549922 493398 549978
rect 492970 532294 493026 532350
rect 493094 532294 493150 532350
rect 493218 532294 493274 532350
rect 493342 532294 493398 532350
rect 492970 532170 493026 532226
rect 493094 532170 493150 532226
rect 493218 532170 493274 532226
rect 493342 532170 493398 532226
rect 492970 532046 493026 532102
rect 493094 532046 493150 532102
rect 493218 532046 493274 532102
rect 493342 532046 493398 532102
rect 492970 531922 493026 531978
rect 493094 531922 493150 531978
rect 493218 531922 493274 531978
rect 493342 531922 493398 531978
rect 507250 597156 507306 597212
rect 507374 597156 507430 597212
rect 507498 597156 507554 597212
rect 507622 597156 507678 597212
rect 507250 597032 507306 597088
rect 507374 597032 507430 597088
rect 507498 597032 507554 597088
rect 507622 597032 507678 597088
rect 507250 596908 507306 596964
rect 507374 596908 507430 596964
rect 507498 596908 507554 596964
rect 507622 596908 507678 596964
rect 507250 596784 507306 596840
rect 507374 596784 507430 596840
rect 507498 596784 507554 596840
rect 507622 596784 507678 596840
rect 507250 580294 507306 580350
rect 507374 580294 507430 580350
rect 507498 580294 507554 580350
rect 507622 580294 507678 580350
rect 507250 580170 507306 580226
rect 507374 580170 507430 580226
rect 507498 580170 507554 580226
rect 507622 580170 507678 580226
rect 507250 580046 507306 580102
rect 507374 580046 507430 580102
rect 507498 580046 507554 580102
rect 507622 580046 507678 580102
rect 507250 579922 507306 579978
rect 507374 579922 507430 579978
rect 507498 579922 507554 579978
rect 507622 579922 507678 579978
rect 507250 562294 507306 562350
rect 507374 562294 507430 562350
rect 507498 562294 507554 562350
rect 507622 562294 507678 562350
rect 507250 562170 507306 562226
rect 507374 562170 507430 562226
rect 507498 562170 507554 562226
rect 507622 562170 507678 562226
rect 507250 562046 507306 562102
rect 507374 562046 507430 562102
rect 507498 562046 507554 562102
rect 507622 562046 507678 562102
rect 507250 561922 507306 561978
rect 507374 561922 507430 561978
rect 507498 561922 507554 561978
rect 507622 561922 507678 561978
rect 507250 544294 507306 544350
rect 507374 544294 507430 544350
rect 507498 544294 507554 544350
rect 507622 544294 507678 544350
rect 507250 544170 507306 544226
rect 507374 544170 507430 544226
rect 507498 544170 507554 544226
rect 507622 544170 507678 544226
rect 507250 544046 507306 544102
rect 507374 544046 507430 544102
rect 507498 544046 507554 544102
rect 507622 544046 507678 544102
rect 507250 543922 507306 543978
rect 507374 543922 507430 543978
rect 507498 543922 507554 543978
rect 507622 543922 507678 543978
rect 507250 526294 507306 526350
rect 507374 526294 507430 526350
rect 507498 526294 507554 526350
rect 507622 526294 507678 526350
rect 507250 526170 507306 526226
rect 507374 526170 507430 526226
rect 507498 526170 507554 526226
rect 507622 526170 507678 526226
rect 507250 526046 507306 526102
rect 507374 526046 507430 526102
rect 507498 526046 507554 526102
rect 507622 526046 507678 526102
rect 507250 525922 507306 525978
rect 507374 525922 507430 525978
rect 507498 525922 507554 525978
rect 507622 525922 507678 525978
rect 510970 598116 511026 598172
rect 511094 598116 511150 598172
rect 511218 598116 511274 598172
rect 511342 598116 511398 598172
rect 510970 597992 511026 598048
rect 511094 597992 511150 598048
rect 511218 597992 511274 598048
rect 511342 597992 511398 598048
rect 510970 597868 511026 597924
rect 511094 597868 511150 597924
rect 511218 597868 511274 597924
rect 511342 597868 511398 597924
rect 510970 597744 511026 597800
rect 511094 597744 511150 597800
rect 511218 597744 511274 597800
rect 511342 597744 511398 597800
rect 510970 586294 511026 586350
rect 511094 586294 511150 586350
rect 511218 586294 511274 586350
rect 511342 586294 511398 586350
rect 510970 586170 511026 586226
rect 511094 586170 511150 586226
rect 511218 586170 511274 586226
rect 511342 586170 511398 586226
rect 510970 586046 511026 586102
rect 511094 586046 511150 586102
rect 511218 586046 511274 586102
rect 511342 586046 511398 586102
rect 510970 585922 511026 585978
rect 511094 585922 511150 585978
rect 511218 585922 511274 585978
rect 511342 585922 511398 585978
rect 510970 568294 511026 568350
rect 511094 568294 511150 568350
rect 511218 568294 511274 568350
rect 511342 568294 511398 568350
rect 510970 568170 511026 568226
rect 511094 568170 511150 568226
rect 511218 568170 511274 568226
rect 511342 568170 511398 568226
rect 510970 568046 511026 568102
rect 511094 568046 511150 568102
rect 511218 568046 511274 568102
rect 511342 568046 511398 568102
rect 510970 567922 511026 567978
rect 511094 567922 511150 567978
rect 511218 567922 511274 567978
rect 511342 567922 511398 567978
rect 510970 550294 511026 550350
rect 511094 550294 511150 550350
rect 511218 550294 511274 550350
rect 511342 550294 511398 550350
rect 510970 550170 511026 550226
rect 511094 550170 511150 550226
rect 511218 550170 511274 550226
rect 511342 550170 511398 550226
rect 510970 550046 511026 550102
rect 511094 550046 511150 550102
rect 511218 550046 511274 550102
rect 511342 550046 511398 550102
rect 510970 549922 511026 549978
rect 511094 549922 511150 549978
rect 511218 549922 511274 549978
rect 511342 549922 511398 549978
rect 510970 532294 511026 532350
rect 511094 532294 511150 532350
rect 511218 532294 511274 532350
rect 511342 532294 511398 532350
rect 510970 532170 511026 532226
rect 511094 532170 511150 532226
rect 511218 532170 511274 532226
rect 511342 532170 511398 532226
rect 510970 532046 511026 532102
rect 511094 532046 511150 532102
rect 511218 532046 511274 532102
rect 511342 532046 511398 532102
rect 510970 531922 511026 531978
rect 511094 531922 511150 531978
rect 511218 531922 511274 531978
rect 511342 531922 511398 531978
rect 525250 597156 525306 597212
rect 525374 597156 525430 597212
rect 525498 597156 525554 597212
rect 525622 597156 525678 597212
rect 525250 597032 525306 597088
rect 525374 597032 525430 597088
rect 525498 597032 525554 597088
rect 525622 597032 525678 597088
rect 525250 596908 525306 596964
rect 525374 596908 525430 596964
rect 525498 596908 525554 596964
rect 525622 596908 525678 596964
rect 525250 596784 525306 596840
rect 525374 596784 525430 596840
rect 525498 596784 525554 596840
rect 525622 596784 525678 596840
rect 525250 580294 525306 580350
rect 525374 580294 525430 580350
rect 525498 580294 525554 580350
rect 525622 580294 525678 580350
rect 525250 580170 525306 580226
rect 525374 580170 525430 580226
rect 525498 580170 525554 580226
rect 525622 580170 525678 580226
rect 525250 580046 525306 580102
rect 525374 580046 525430 580102
rect 525498 580046 525554 580102
rect 525622 580046 525678 580102
rect 525250 579922 525306 579978
rect 525374 579922 525430 579978
rect 525498 579922 525554 579978
rect 525622 579922 525678 579978
rect 525250 562294 525306 562350
rect 525374 562294 525430 562350
rect 525498 562294 525554 562350
rect 525622 562294 525678 562350
rect 525250 562170 525306 562226
rect 525374 562170 525430 562226
rect 525498 562170 525554 562226
rect 525622 562170 525678 562226
rect 525250 562046 525306 562102
rect 525374 562046 525430 562102
rect 525498 562046 525554 562102
rect 525622 562046 525678 562102
rect 525250 561922 525306 561978
rect 525374 561922 525430 561978
rect 525498 561922 525554 561978
rect 525622 561922 525678 561978
rect 525250 544294 525306 544350
rect 525374 544294 525430 544350
rect 525498 544294 525554 544350
rect 525622 544294 525678 544350
rect 525250 544170 525306 544226
rect 525374 544170 525430 544226
rect 525498 544170 525554 544226
rect 525622 544170 525678 544226
rect 525250 544046 525306 544102
rect 525374 544046 525430 544102
rect 525498 544046 525554 544102
rect 525622 544046 525678 544102
rect 525250 543922 525306 543978
rect 525374 543922 525430 543978
rect 525498 543922 525554 543978
rect 525622 543922 525678 543978
rect 525250 526294 525306 526350
rect 525374 526294 525430 526350
rect 525498 526294 525554 526350
rect 525622 526294 525678 526350
rect 525250 526170 525306 526226
rect 525374 526170 525430 526226
rect 525498 526170 525554 526226
rect 525622 526170 525678 526226
rect 525250 526046 525306 526102
rect 525374 526046 525430 526102
rect 525498 526046 525554 526102
rect 525622 526046 525678 526102
rect 525250 525922 525306 525978
rect 525374 525922 525430 525978
rect 525498 525922 525554 525978
rect 525622 525922 525678 525978
rect 6970 514294 7026 514350
rect 7094 514294 7150 514350
rect 7218 514294 7274 514350
rect 7342 514294 7398 514350
rect 6970 514170 7026 514226
rect 7094 514170 7150 514226
rect 7218 514170 7274 514226
rect 7342 514170 7398 514226
rect 6970 514046 7026 514102
rect 7094 514046 7150 514102
rect 7218 514046 7274 514102
rect 7342 514046 7398 514102
rect 6970 513922 7026 513978
rect 7094 513922 7150 513978
rect 7218 513922 7274 513978
rect 7342 513922 7398 513978
rect 39878 514294 39934 514350
rect 40002 514294 40058 514350
rect 39878 514170 39934 514226
rect 40002 514170 40058 514226
rect 39878 514046 39934 514102
rect 40002 514046 40058 514102
rect 39878 513922 39934 513978
rect 40002 513922 40058 513978
rect 70598 514294 70654 514350
rect 70722 514294 70778 514350
rect 70598 514170 70654 514226
rect 70722 514170 70778 514226
rect 70598 514046 70654 514102
rect 70722 514046 70778 514102
rect 70598 513922 70654 513978
rect 70722 513922 70778 513978
rect 101318 514294 101374 514350
rect 101442 514294 101498 514350
rect 101318 514170 101374 514226
rect 101442 514170 101498 514226
rect 101318 514046 101374 514102
rect 101442 514046 101498 514102
rect 101318 513922 101374 513978
rect 101442 513922 101498 513978
rect 132038 514294 132094 514350
rect 132162 514294 132218 514350
rect 132038 514170 132094 514226
rect 132162 514170 132218 514226
rect 132038 514046 132094 514102
rect 132162 514046 132218 514102
rect 132038 513922 132094 513978
rect 132162 513922 132218 513978
rect 162758 514294 162814 514350
rect 162882 514294 162938 514350
rect 162758 514170 162814 514226
rect 162882 514170 162938 514226
rect 162758 514046 162814 514102
rect 162882 514046 162938 514102
rect 162758 513922 162814 513978
rect 162882 513922 162938 513978
rect 193478 514294 193534 514350
rect 193602 514294 193658 514350
rect 193478 514170 193534 514226
rect 193602 514170 193658 514226
rect 193478 514046 193534 514102
rect 193602 514046 193658 514102
rect 193478 513922 193534 513978
rect 193602 513922 193658 513978
rect 224198 514294 224254 514350
rect 224322 514294 224378 514350
rect 224198 514170 224254 514226
rect 224322 514170 224378 514226
rect 224198 514046 224254 514102
rect 224322 514046 224378 514102
rect 224198 513922 224254 513978
rect 224322 513922 224378 513978
rect 254918 514294 254974 514350
rect 255042 514294 255098 514350
rect 254918 514170 254974 514226
rect 255042 514170 255098 514226
rect 254918 514046 254974 514102
rect 255042 514046 255098 514102
rect 254918 513922 254974 513978
rect 255042 513922 255098 513978
rect 285638 514294 285694 514350
rect 285762 514294 285818 514350
rect 285638 514170 285694 514226
rect 285762 514170 285818 514226
rect 285638 514046 285694 514102
rect 285762 514046 285818 514102
rect 285638 513922 285694 513978
rect 285762 513922 285818 513978
rect 316358 514294 316414 514350
rect 316482 514294 316538 514350
rect 316358 514170 316414 514226
rect 316482 514170 316538 514226
rect 316358 514046 316414 514102
rect 316482 514046 316538 514102
rect 316358 513922 316414 513978
rect 316482 513922 316538 513978
rect 347078 514294 347134 514350
rect 347202 514294 347258 514350
rect 347078 514170 347134 514226
rect 347202 514170 347258 514226
rect 347078 514046 347134 514102
rect 347202 514046 347258 514102
rect 347078 513922 347134 513978
rect 347202 513922 347258 513978
rect 377798 514294 377854 514350
rect 377922 514294 377978 514350
rect 377798 514170 377854 514226
rect 377922 514170 377978 514226
rect 377798 514046 377854 514102
rect 377922 514046 377978 514102
rect 377798 513922 377854 513978
rect 377922 513922 377978 513978
rect 408518 514294 408574 514350
rect 408642 514294 408698 514350
rect 408518 514170 408574 514226
rect 408642 514170 408698 514226
rect 408518 514046 408574 514102
rect 408642 514046 408698 514102
rect 408518 513922 408574 513978
rect 408642 513922 408698 513978
rect 439238 514294 439294 514350
rect 439362 514294 439418 514350
rect 439238 514170 439294 514226
rect 439362 514170 439418 514226
rect 439238 514046 439294 514102
rect 439362 514046 439418 514102
rect 439238 513922 439294 513978
rect 439362 513922 439418 513978
rect 469958 514294 470014 514350
rect 470082 514294 470138 514350
rect 469958 514170 470014 514226
rect 470082 514170 470138 514226
rect 469958 514046 470014 514102
rect 470082 514046 470138 514102
rect 469958 513922 470014 513978
rect 470082 513922 470138 513978
rect 500678 514294 500734 514350
rect 500802 514294 500858 514350
rect 500678 514170 500734 514226
rect 500802 514170 500858 514226
rect 500678 514046 500734 514102
rect 500802 514046 500858 514102
rect 500678 513922 500734 513978
rect 500802 513922 500858 513978
rect 24518 508294 24574 508350
rect 24642 508294 24698 508350
rect 24518 508170 24574 508226
rect 24642 508170 24698 508226
rect 24518 508046 24574 508102
rect 24642 508046 24698 508102
rect 24518 507922 24574 507978
rect 24642 507922 24698 507978
rect 55238 508294 55294 508350
rect 55362 508294 55418 508350
rect 55238 508170 55294 508226
rect 55362 508170 55418 508226
rect 55238 508046 55294 508102
rect 55362 508046 55418 508102
rect 55238 507922 55294 507978
rect 55362 507922 55418 507978
rect 85958 508294 86014 508350
rect 86082 508294 86138 508350
rect 85958 508170 86014 508226
rect 86082 508170 86138 508226
rect 85958 508046 86014 508102
rect 86082 508046 86138 508102
rect 85958 507922 86014 507978
rect 86082 507922 86138 507978
rect 116678 508294 116734 508350
rect 116802 508294 116858 508350
rect 116678 508170 116734 508226
rect 116802 508170 116858 508226
rect 116678 508046 116734 508102
rect 116802 508046 116858 508102
rect 116678 507922 116734 507978
rect 116802 507922 116858 507978
rect 147398 508294 147454 508350
rect 147522 508294 147578 508350
rect 147398 508170 147454 508226
rect 147522 508170 147578 508226
rect 147398 508046 147454 508102
rect 147522 508046 147578 508102
rect 147398 507922 147454 507978
rect 147522 507922 147578 507978
rect 178118 508294 178174 508350
rect 178242 508294 178298 508350
rect 178118 508170 178174 508226
rect 178242 508170 178298 508226
rect 178118 508046 178174 508102
rect 178242 508046 178298 508102
rect 178118 507922 178174 507978
rect 178242 507922 178298 507978
rect 208838 508294 208894 508350
rect 208962 508294 209018 508350
rect 208838 508170 208894 508226
rect 208962 508170 209018 508226
rect 208838 508046 208894 508102
rect 208962 508046 209018 508102
rect 208838 507922 208894 507978
rect 208962 507922 209018 507978
rect 239558 508294 239614 508350
rect 239682 508294 239738 508350
rect 239558 508170 239614 508226
rect 239682 508170 239738 508226
rect 239558 508046 239614 508102
rect 239682 508046 239738 508102
rect 239558 507922 239614 507978
rect 239682 507922 239738 507978
rect 270278 508294 270334 508350
rect 270402 508294 270458 508350
rect 270278 508170 270334 508226
rect 270402 508170 270458 508226
rect 270278 508046 270334 508102
rect 270402 508046 270458 508102
rect 270278 507922 270334 507978
rect 270402 507922 270458 507978
rect 300998 508294 301054 508350
rect 301122 508294 301178 508350
rect 300998 508170 301054 508226
rect 301122 508170 301178 508226
rect 300998 508046 301054 508102
rect 301122 508046 301178 508102
rect 300998 507922 301054 507978
rect 301122 507922 301178 507978
rect 331718 508294 331774 508350
rect 331842 508294 331898 508350
rect 331718 508170 331774 508226
rect 331842 508170 331898 508226
rect 331718 508046 331774 508102
rect 331842 508046 331898 508102
rect 331718 507922 331774 507978
rect 331842 507922 331898 507978
rect 362438 508294 362494 508350
rect 362562 508294 362618 508350
rect 362438 508170 362494 508226
rect 362562 508170 362618 508226
rect 362438 508046 362494 508102
rect 362562 508046 362618 508102
rect 362438 507922 362494 507978
rect 362562 507922 362618 507978
rect 393158 508294 393214 508350
rect 393282 508294 393338 508350
rect 393158 508170 393214 508226
rect 393282 508170 393338 508226
rect 393158 508046 393214 508102
rect 393282 508046 393338 508102
rect 393158 507922 393214 507978
rect 393282 507922 393338 507978
rect 423878 508294 423934 508350
rect 424002 508294 424058 508350
rect 423878 508170 423934 508226
rect 424002 508170 424058 508226
rect 423878 508046 423934 508102
rect 424002 508046 424058 508102
rect 423878 507922 423934 507978
rect 424002 507922 424058 507978
rect 454598 508294 454654 508350
rect 454722 508294 454778 508350
rect 454598 508170 454654 508226
rect 454722 508170 454778 508226
rect 454598 508046 454654 508102
rect 454722 508046 454778 508102
rect 454598 507922 454654 507978
rect 454722 507922 454778 507978
rect 485318 508294 485374 508350
rect 485442 508294 485498 508350
rect 485318 508170 485374 508226
rect 485442 508170 485498 508226
rect 485318 508046 485374 508102
rect 485442 508046 485498 508102
rect 485318 507922 485374 507978
rect 485442 507922 485498 507978
rect 516038 508294 516094 508350
rect 516162 508294 516218 508350
rect 516038 508170 516094 508226
rect 516162 508170 516218 508226
rect 516038 508046 516094 508102
rect 516162 508046 516218 508102
rect 516038 507922 516094 507978
rect 516162 507922 516218 507978
rect 525250 508294 525306 508350
rect 525374 508294 525430 508350
rect 525498 508294 525554 508350
rect 525622 508294 525678 508350
rect 525250 508170 525306 508226
rect 525374 508170 525430 508226
rect 525498 508170 525554 508226
rect 525622 508170 525678 508226
rect 525250 508046 525306 508102
rect 525374 508046 525430 508102
rect 525498 508046 525554 508102
rect 525622 508046 525678 508102
rect 525250 507922 525306 507978
rect 525374 507922 525430 507978
rect 525498 507922 525554 507978
rect 525622 507922 525678 507978
rect 6970 496294 7026 496350
rect 7094 496294 7150 496350
rect 7218 496294 7274 496350
rect 7342 496294 7398 496350
rect 6970 496170 7026 496226
rect 7094 496170 7150 496226
rect 7218 496170 7274 496226
rect 7342 496170 7398 496226
rect 6970 496046 7026 496102
rect 7094 496046 7150 496102
rect 7218 496046 7274 496102
rect 7342 496046 7398 496102
rect 6970 495922 7026 495978
rect 7094 495922 7150 495978
rect 7218 495922 7274 495978
rect 7342 495922 7398 495978
rect 39878 496294 39934 496350
rect 40002 496294 40058 496350
rect 39878 496170 39934 496226
rect 40002 496170 40058 496226
rect 39878 496046 39934 496102
rect 40002 496046 40058 496102
rect 39878 495922 39934 495978
rect 40002 495922 40058 495978
rect 70598 496294 70654 496350
rect 70722 496294 70778 496350
rect 70598 496170 70654 496226
rect 70722 496170 70778 496226
rect 70598 496046 70654 496102
rect 70722 496046 70778 496102
rect 70598 495922 70654 495978
rect 70722 495922 70778 495978
rect 101318 496294 101374 496350
rect 101442 496294 101498 496350
rect 101318 496170 101374 496226
rect 101442 496170 101498 496226
rect 101318 496046 101374 496102
rect 101442 496046 101498 496102
rect 101318 495922 101374 495978
rect 101442 495922 101498 495978
rect 132038 496294 132094 496350
rect 132162 496294 132218 496350
rect 132038 496170 132094 496226
rect 132162 496170 132218 496226
rect 132038 496046 132094 496102
rect 132162 496046 132218 496102
rect 132038 495922 132094 495978
rect 132162 495922 132218 495978
rect 162758 496294 162814 496350
rect 162882 496294 162938 496350
rect 162758 496170 162814 496226
rect 162882 496170 162938 496226
rect 162758 496046 162814 496102
rect 162882 496046 162938 496102
rect 162758 495922 162814 495978
rect 162882 495922 162938 495978
rect 193478 496294 193534 496350
rect 193602 496294 193658 496350
rect 193478 496170 193534 496226
rect 193602 496170 193658 496226
rect 193478 496046 193534 496102
rect 193602 496046 193658 496102
rect 193478 495922 193534 495978
rect 193602 495922 193658 495978
rect 224198 496294 224254 496350
rect 224322 496294 224378 496350
rect 224198 496170 224254 496226
rect 224322 496170 224378 496226
rect 224198 496046 224254 496102
rect 224322 496046 224378 496102
rect 224198 495922 224254 495978
rect 224322 495922 224378 495978
rect 254918 496294 254974 496350
rect 255042 496294 255098 496350
rect 254918 496170 254974 496226
rect 255042 496170 255098 496226
rect 254918 496046 254974 496102
rect 255042 496046 255098 496102
rect 254918 495922 254974 495978
rect 255042 495922 255098 495978
rect 285638 496294 285694 496350
rect 285762 496294 285818 496350
rect 285638 496170 285694 496226
rect 285762 496170 285818 496226
rect 285638 496046 285694 496102
rect 285762 496046 285818 496102
rect 285638 495922 285694 495978
rect 285762 495922 285818 495978
rect 316358 496294 316414 496350
rect 316482 496294 316538 496350
rect 316358 496170 316414 496226
rect 316482 496170 316538 496226
rect 316358 496046 316414 496102
rect 316482 496046 316538 496102
rect 316358 495922 316414 495978
rect 316482 495922 316538 495978
rect 347078 496294 347134 496350
rect 347202 496294 347258 496350
rect 347078 496170 347134 496226
rect 347202 496170 347258 496226
rect 347078 496046 347134 496102
rect 347202 496046 347258 496102
rect 347078 495922 347134 495978
rect 347202 495922 347258 495978
rect 377798 496294 377854 496350
rect 377922 496294 377978 496350
rect 377798 496170 377854 496226
rect 377922 496170 377978 496226
rect 377798 496046 377854 496102
rect 377922 496046 377978 496102
rect 377798 495922 377854 495978
rect 377922 495922 377978 495978
rect 408518 496294 408574 496350
rect 408642 496294 408698 496350
rect 408518 496170 408574 496226
rect 408642 496170 408698 496226
rect 408518 496046 408574 496102
rect 408642 496046 408698 496102
rect 408518 495922 408574 495978
rect 408642 495922 408698 495978
rect 439238 496294 439294 496350
rect 439362 496294 439418 496350
rect 439238 496170 439294 496226
rect 439362 496170 439418 496226
rect 439238 496046 439294 496102
rect 439362 496046 439418 496102
rect 439238 495922 439294 495978
rect 439362 495922 439418 495978
rect 469958 496294 470014 496350
rect 470082 496294 470138 496350
rect 469958 496170 470014 496226
rect 470082 496170 470138 496226
rect 469958 496046 470014 496102
rect 470082 496046 470138 496102
rect 469958 495922 470014 495978
rect 470082 495922 470138 495978
rect 500678 496294 500734 496350
rect 500802 496294 500858 496350
rect 500678 496170 500734 496226
rect 500802 496170 500858 496226
rect 500678 496046 500734 496102
rect 500802 496046 500858 496102
rect 500678 495922 500734 495978
rect 500802 495922 500858 495978
rect 24518 490294 24574 490350
rect 24642 490294 24698 490350
rect 24518 490170 24574 490226
rect 24642 490170 24698 490226
rect 24518 490046 24574 490102
rect 24642 490046 24698 490102
rect 24518 489922 24574 489978
rect 24642 489922 24698 489978
rect 55238 490294 55294 490350
rect 55362 490294 55418 490350
rect 55238 490170 55294 490226
rect 55362 490170 55418 490226
rect 55238 490046 55294 490102
rect 55362 490046 55418 490102
rect 55238 489922 55294 489978
rect 55362 489922 55418 489978
rect 85958 490294 86014 490350
rect 86082 490294 86138 490350
rect 85958 490170 86014 490226
rect 86082 490170 86138 490226
rect 85958 490046 86014 490102
rect 86082 490046 86138 490102
rect 85958 489922 86014 489978
rect 86082 489922 86138 489978
rect 116678 490294 116734 490350
rect 116802 490294 116858 490350
rect 116678 490170 116734 490226
rect 116802 490170 116858 490226
rect 116678 490046 116734 490102
rect 116802 490046 116858 490102
rect 116678 489922 116734 489978
rect 116802 489922 116858 489978
rect 147398 490294 147454 490350
rect 147522 490294 147578 490350
rect 147398 490170 147454 490226
rect 147522 490170 147578 490226
rect 147398 490046 147454 490102
rect 147522 490046 147578 490102
rect 147398 489922 147454 489978
rect 147522 489922 147578 489978
rect 178118 490294 178174 490350
rect 178242 490294 178298 490350
rect 178118 490170 178174 490226
rect 178242 490170 178298 490226
rect 178118 490046 178174 490102
rect 178242 490046 178298 490102
rect 178118 489922 178174 489978
rect 178242 489922 178298 489978
rect 208838 490294 208894 490350
rect 208962 490294 209018 490350
rect 208838 490170 208894 490226
rect 208962 490170 209018 490226
rect 208838 490046 208894 490102
rect 208962 490046 209018 490102
rect 208838 489922 208894 489978
rect 208962 489922 209018 489978
rect 239558 490294 239614 490350
rect 239682 490294 239738 490350
rect 239558 490170 239614 490226
rect 239682 490170 239738 490226
rect 239558 490046 239614 490102
rect 239682 490046 239738 490102
rect 239558 489922 239614 489978
rect 239682 489922 239738 489978
rect 270278 490294 270334 490350
rect 270402 490294 270458 490350
rect 270278 490170 270334 490226
rect 270402 490170 270458 490226
rect 270278 490046 270334 490102
rect 270402 490046 270458 490102
rect 270278 489922 270334 489978
rect 270402 489922 270458 489978
rect 300998 490294 301054 490350
rect 301122 490294 301178 490350
rect 300998 490170 301054 490226
rect 301122 490170 301178 490226
rect 300998 490046 301054 490102
rect 301122 490046 301178 490102
rect 300998 489922 301054 489978
rect 301122 489922 301178 489978
rect 331718 490294 331774 490350
rect 331842 490294 331898 490350
rect 331718 490170 331774 490226
rect 331842 490170 331898 490226
rect 331718 490046 331774 490102
rect 331842 490046 331898 490102
rect 331718 489922 331774 489978
rect 331842 489922 331898 489978
rect 362438 490294 362494 490350
rect 362562 490294 362618 490350
rect 362438 490170 362494 490226
rect 362562 490170 362618 490226
rect 362438 490046 362494 490102
rect 362562 490046 362618 490102
rect 362438 489922 362494 489978
rect 362562 489922 362618 489978
rect 393158 490294 393214 490350
rect 393282 490294 393338 490350
rect 393158 490170 393214 490226
rect 393282 490170 393338 490226
rect 393158 490046 393214 490102
rect 393282 490046 393338 490102
rect 393158 489922 393214 489978
rect 393282 489922 393338 489978
rect 423878 490294 423934 490350
rect 424002 490294 424058 490350
rect 423878 490170 423934 490226
rect 424002 490170 424058 490226
rect 423878 490046 423934 490102
rect 424002 490046 424058 490102
rect 423878 489922 423934 489978
rect 424002 489922 424058 489978
rect 454598 490294 454654 490350
rect 454722 490294 454778 490350
rect 454598 490170 454654 490226
rect 454722 490170 454778 490226
rect 454598 490046 454654 490102
rect 454722 490046 454778 490102
rect 454598 489922 454654 489978
rect 454722 489922 454778 489978
rect 485318 490294 485374 490350
rect 485442 490294 485498 490350
rect 485318 490170 485374 490226
rect 485442 490170 485498 490226
rect 485318 490046 485374 490102
rect 485442 490046 485498 490102
rect 485318 489922 485374 489978
rect 485442 489922 485498 489978
rect 516038 490294 516094 490350
rect 516162 490294 516218 490350
rect 516038 490170 516094 490226
rect 516162 490170 516218 490226
rect 516038 490046 516094 490102
rect 516162 490046 516218 490102
rect 516038 489922 516094 489978
rect 516162 489922 516218 489978
rect 525250 490294 525306 490350
rect 525374 490294 525430 490350
rect 525498 490294 525554 490350
rect 525622 490294 525678 490350
rect 525250 490170 525306 490226
rect 525374 490170 525430 490226
rect 525498 490170 525554 490226
rect 525622 490170 525678 490226
rect 525250 490046 525306 490102
rect 525374 490046 525430 490102
rect 525498 490046 525554 490102
rect 525622 490046 525678 490102
rect 525250 489922 525306 489978
rect 525374 489922 525430 489978
rect 525498 489922 525554 489978
rect 525622 489922 525678 489978
rect 6970 478294 7026 478350
rect 7094 478294 7150 478350
rect 7218 478294 7274 478350
rect 7342 478294 7398 478350
rect 6970 478170 7026 478226
rect 7094 478170 7150 478226
rect 7218 478170 7274 478226
rect 7342 478170 7398 478226
rect 6970 478046 7026 478102
rect 7094 478046 7150 478102
rect 7218 478046 7274 478102
rect 7342 478046 7398 478102
rect 6970 477922 7026 477978
rect 7094 477922 7150 477978
rect 7218 477922 7274 477978
rect 7342 477922 7398 477978
rect 39878 478294 39934 478350
rect 40002 478294 40058 478350
rect 39878 478170 39934 478226
rect 40002 478170 40058 478226
rect 39878 478046 39934 478102
rect 40002 478046 40058 478102
rect 39878 477922 39934 477978
rect 40002 477922 40058 477978
rect 70598 478294 70654 478350
rect 70722 478294 70778 478350
rect 70598 478170 70654 478226
rect 70722 478170 70778 478226
rect 70598 478046 70654 478102
rect 70722 478046 70778 478102
rect 70598 477922 70654 477978
rect 70722 477922 70778 477978
rect 101318 478294 101374 478350
rect 101442 478294 101498 478350
rect 101318 478170 101374 478226
rect 101442 478170 101498 478226
rect 101318 478046 101374 478102
rect 101442 478046 101498 478102
rect 101318 477922 101374 477978
rect 101442 477922 101498 477978
rect 132038 478294 132094 478350
rect 132162 478294 132218 478350
rect 132038 478170 132094 478226
rect 132162 478170 132218 478226
rect 132038 478046 132094 478102
rect 132162 478046 132218 478102
rect 132038 477922 132094 477978
rect 132162 477922 132218 477978
rect 162758 478294 162814 478350
rect 162882 478294 162938 478350
rect 162758 478170 162814 478226
rect 162882 478170 162938 478226
rect 162758 478046 162814 478102
rect 162882 478046 162938 478102
rect 162758 477922 162814 477978
rect 162882 477922 162938 477978
rect 193478 478294 193534 478350
rect 193602 478294 193658 478350
rect 193478 478170 193534 478226
rect 193602 478170 193658 478226
rect 193478 478046 193534 478102
rect 193602 478046 193658 478102
rect 193478 477922 193534 477978
rect 193602 477922 193658 477978
rect 224198 478294 224254 478350
rect 224322 478294 224378 478350
rect 224198 478170 224254 478226
rect 224322 478170 224378 478226
rect 224198 478046 224254 478102
rect 224322 478046 224378 478102
rect 224198 477922 224254 477978
rect 224322 477922 224378 477978
rect 254918 478294 254974 478350
rect 255042 478294 255098 478350
rect 254918 478170 254974 478226
rect 255042 478170 255098 478226
rect 254918 478046 254974 478102
rect 255042 478046 255098 478102
rect 254918 477922 254974 477978
rect 255042 477922 255098 477978
rect 285638 478294 285694 478350
rect 285762 478294 285818 478350
rect 285638 478170 285694 478226
rect 285762 478170 285818 478226
rect 285638 478046 285694 478102
rect 285762 478046 285818 478102
rect 285638 477922 285694 477978
rect 285762 477922 285818 477978
rect 316358 478294 316414 478350
rect 316482 478294 316538 478350
rect 316358 478170 316414 478226
rect 316482 478170 316538 478226
rect 316358 478046 316414 478102
rect 316482 478046 316538 478102
rect 316358 477922 316414 477978
rect 316482 477922 316538 477978
rect 347078 478294 347134 478350
rect 347202 478294 347258 478350
rect 347078 478170 347134 478226
rect 347202 478170 347258 478226
rect 347078 478046 347134 478102
rect 347202 478046 347258 478102
rect 347078 477922 347134 477978
rect 347202 477922 347258 477978
rect 377798 478294 377854 478350
rect 377922 478294 377978 478350
rect 377798 478170 377854 478226
rect 377922 478170 377978 478226
rect 377798 478046 377854 478102
rect 377922 478046 377978 478102
rect 377798 477922 377854 477978
rect 377922 477922 377978 477978
rect 408518 478294 408574 478350
rect 408642 478294 408698 478350
rect 408518 478170 408574 478226
rect 408642 478170 408698 478226
rect 408518 478046 408574 478102
rect 408642 478046 408698 478102
rect 408518 477922 408574 477978
rect 408642 477922 408698 477978
rect 439238 478294 439294 478350
rect 439362 478294 439418 478350
rect 439238 478170 439294 478226
rect 439362 478170 439418 478226
rect 439238 478046 439294 478102
rect 439362 478046 439418 478102
rect 439238 477922 439294 477978
rect 439362 477922 439418 477978
rect 469958 478294 470014 478350
rect 470082 478294 470138 478350
rect 469958 478170 470014 478226
rect 470082 478170 470138 478226
rect 469958 478046 470014 478102
rect 470082 478046 470138 478102
rect 469958 477922 470014 477978
rect 470082 477922 470138 477978
rect 500678 478294 500734 478350
rect 500802 478294 500858 478350
rect 500678 478170 500734 478226
rect 500802 478170 500858 478226
rect 500678 478046 500734 478102
rect 500802 478046 500858 478102
rect 500678 477922 500734 477978
rect 500802 477922 500858 477978
rect 24518 472294 24574 472350
rect 24642 472294 24698 472350
rect 24518 472170 24574 472226
rect 24642 472170 24698 472226
rect 24518 472046 24574 472102
rect 24642 472046 24698 472102
rect 24518 471922 24574 471978
rect 24642 471922 24698 471978
rect 55238 472294 55294 472350
rect 55362 472294 55418 472350
rect 55238 472170 55294 472226
rect 55362 472170 55418 472226
rect 55238 472046 55294 472102
rect 55362 472046 55418 472102
rect 55238 471922 55294 471978
rect 55362 471922 55418 471978
rect 85958 472294 86014 472350
rect 86082 472294 86138 472350
rect 85958 472170 86014 472226
rect 86082 472170 86138 472226
rect 85958 472046 86014 472102
rect 86082 472046 86138 472102
rect 85958 471922 86014 471978
rect 86082 471922 86138 471978
rect 116678 472294 116734 472350
rect 116802 472294 116858 472350
rect 116678 472170 116734 472226
rect 116802 472170 116858 472226
rect 116678 472046 116734 472102
rect 116802 472046 116858 472102
rect 116678 471922 116734 471978
rect 116802 471922 116858 471978
rect 147398 472294 147454 472350
rect 147522 472294 147578 472350
rect 147398 472170 147454 472226
rect 147522 472170 147578 472226
rect 147398 472046 147454 472102
rect 147522 472046 147578 472102
rect 147398 471922 147454 471978
rect 147522 471922 147578 471978
rect 178118 472294 178174 472350
rect 178242 472294 178298 472350
rect 178118 472170 178174 472226
rect 178242 472170 178298 472226
rect 178118 472046 178174 472102
rect 178242 472046 178298 472102
rect 178118 471922 178174 471978
rect 178242 471922 178298 471978
rect 208838 472294 208894 472350
rect 208962 472294 209018 472350
rect 208838 472170 208894 472226
rect 208962 472170 209018 472226
rect 208838 472046 208894 472102
rect 208962 472046 209018 472102
rect 208838 471922 208894 471978
rect 208962 471922 209018 471978
rect 239558 472294 239614 472350
rect 239682 472294 239738 472350
rect 239558 472170 239614 472226
rect 239682 472170 239738 472226
rect 239558 472046 239614 472102
rect 239682 472046 239738 472102
rect 239558 471922 239614 471978
rect 239682 471922 239738 471978
rect 270278 472294 270334 472350
rect 270402 472294 270458 472350
rect 270278 472170 270334 472226
rect 270402 472170 270458 472226
rect 270278 472046 270334 472102
rect 270402 472046 270458 472102
rect 270278 471922 270334 471978
rect 270402 471922 270458 471978
rect 300998 472294 301054 472350
rect 301122 472294 301178 472350
rect 300998 472170 301054 472226
rect 301122 472170 301178 472226
rect 300998 472046 301054 472102
rect 301122 472046 301178 472102
rect 300998 471922 301054 471978
rect 301122 471922 301178 471978
rect 331718 472294 331774 472350
rect 331842 472294 331898 472350
rect 331718 472170 331774 472226
rect 331842 472170 331898 472226
rect 331718 472046 331774 472102
rect 331842 472046 331898 472102
rect 331718 471922 331774 471978
rect 331842 471922 331898 471978
rect 362438 472294 362494 472350
rect 362562 472294 362618 472350
rect 362438 472170 362494 472226
rect 362562 472170 362618 472226
rect 362438 472046 362494 472102
rect 362562 472046 362618 472102
rect 362438 471922 362494 471978
rect 362562 471922 362618 471978
rect 393158 472294 393214 472350
rect 393282 472294 393338 472350
rect 393158 472170 393214 472226
rect 393282 472170 393338 472226
rect 393158 472046 393214 472102
rect 393282 472046 393338 472102
rect 393158 471922 393214 471978
rect 393282 471922 393338 471978
rect 423878 472294 423934 472350
rect 424002 472294 424058 472350
rect 423878 472170 423934 472226
rect 424002 472170 424058 472226
rect 423878 472046 423934 472102
rect 424002 472046 424058 472102
rect 423878 471922 423934 471978
rect 424002 471922 424058 471978
rect 454598 472294 454654 472350
rect 454722 472294 454778 472350
rect 454598 472170 454654 472226
rect 454722 472170 454778 472226
rect 454598 472046 454654 472102
rect 454722 472046 454778 472102
rect 454598 471922 454654 471978
rect 454722 471922 454778 471978
rect 485318 472294 485374 472350
rect 485442 472294 485498 472350
rect 485318 472170 485374 472226
rect 485442 472170 485498 472226
rect 485318 472046 485374 472102
rect 485442 472046 485498 472102
rect 485318 471922 485374 471978
rect 485442 471922 485498 471978
rect 516038 472294 516094 472350
rect 516162 472294 516218 472350
rect 516038 472170 516094 472226
rect 516162 472170 516218 472226
rect 516038 472046 516094 472102
rect 516162 472046 516218 472102
rect 516038 471922 516094 471978
rect 516162 471922 516218 471978
rect 525250 472294 525306 472350
rect 525374 472294 525430 472350
rect 525498 472294 525554 472350
rect 525622 472294 525678 472350
rect 525250 472170 525306 472226
rect 525374 472170 525430 472226
rect 525498 472170 525554 472226
rect 525622 472170 525678 472226
rect 525250 472046 525306 472102
rect 525374 472046 525430 472102
rect 525498 472046 525554 472102
rect 525622 472046 525678 472102
rect 525250 471922 525306 471978
rect 525374 471922 525430 471978
rect 525498 471922 525554 471978
rect 525622 471922 525678 471978
rect 6970 460294 7026 460350
rect 7094 460294 7150 460350
rect 7218 460294 7274 460350
rect 7342 460294 7398 460350
rect 6970 460170 7026 460226
rect 7094 460170 7150 460226
rect 7218 460170 7274 460226
rect 7342 460170 7398 460226
rect 6970 460046 7026 460102
rect 7094 460046 7150 460102
rect 7218 460046 7274 460102
rect 7342 460046 7398 460102
rect 6970 459922 7026 459978
rect 7094 459922 7150 459978
rect 7218 459922 7274 459978
rect 7342 459922 7398 459978
rect 39878 460294 39934 460350
rect 40002 460294 40058 460350
rect 39878 460170 39934 460226
rect 40002 460170 40058 460226
rect 39878 460046 39934 460102
rect 40002 460046 40058 460102
rect 39878 459922 39934 459978
rect 40002 459922 40058 459978
rect 70598 460294 70654 460350
rect 70722 460294 70778 460350
rect 70598 460170 70654 460226
rect 70722 460170 70778 460226
rect 70598 460046 70654 460102
rect 70722 460046 70778 460102
rect 70598 459922 70654 459978
rect 70722 459922 70778 459978
rect 101318 460294 101374 460350
rect 101442 460294 101498 460350
rect 101318 460170 101374 460226
rect 101442 460170 101498 460226
rect 101318 460046 101374 460102
rect 101442 460046 101498 460102
rect 101318 459922 101374 459978
rect 101442 459922 101498 459978
rect 132038 460294 132094 460350
rect 132162 460294 132218 460350
rect 132038 460170 132094 460226
rect 132162 460170 132218 460226
rect 132038 460046 132094 460102
rect 132162 460046 132218 460102
rect 132038 459922 132094 459978
rect 132162 459922 132218 459978
rect 162758 460294 162814 460350
rect 162882 460294 162938 460350
rect 162758 460170 162814 460226
rect 162882 460170 162938 460226
rect 162758 460046 162814 460102
rect 162882 460046 162938 460102
rect 162758 459922 162814 459978
rect 162882 459922 162938 459978
rect 193478 460294 193534 460350
rect 193602 460294 193658 460350
rect 193478 460170 193534 460226
rect 193602 460170 193658 460226
rect 193478 460046 193534 460102
rect 193602 460046 193658 460102
rect 193478 459922 193534 459978
rect 193602 459922 193658 459978
rect 224198 460294 224254 460350
rect 224322 460294 224378 460350
rect 224198 460170 224254 460226
rect 224322 460170 224378 460226
rect 224198 460046 224254 460102
rect 224322 460046 224378 460102
rect 224198 459922 224254 459978
rect 224322 459922 224378 459978
rect 254918 460294 254974 460350
rect 255042 460294 255098 460350
rect 254918 460170 254974 460226
rect 255042 460170 255098 460226
rect 254918 460046 254974 460102
rect 255042 460046 255098 460102
rect 254918 459922 254974 459978
rect 255042 459922 255098 459978
rect 285638 460294 285694 460350
rect 285762 460294 285818 460350
rect 285638 460170 285694 460226
rect 285762 460170 285818 460226
rect 285638 460046 285694 460102
rect 285762 460046 285818 460102
rect 285638 459922 285694 459978
rect 285762 459922 285818 459978
rect 316358 460294 316414 460350
rect 316482 460294 316538 460350
rect 316358 460170 316414 460226
rect 316482 460170 316538 460226
rect 316358 460046 316414 460102
rect 316482 460046 316538 460102
rect 316358 459922 316414 459978
rect 316482 459922 316538 459978
rect 347078 460294 347134 460350
rect 347202 460294 347258 460350
rect 347078 460170 347134 460226
rect 347202 460170 347258 460226
rect 347078 460046 347134 460102
rect 347202 460046 347258 460102
rect 347078 459922 347134 459978
rect 347202 459922 347258 459978
rect 377798 460294 377854 460350
rect 377922 460294 377978 460350
rect 377798 460170 377854 460226
rect 377922 460170 377978 460226
rect 377798 460046 377854 460102
rect 377922 460046 377978 460102
rect 377798 459922 377854 459978
rect 377922 459922 377978 459978
rect 408518 460294 408574 460350
rect 408642 460294 408698 460350
rect 408518 460170 408574 460226
rect 408642 460170 408698 460226
rect 408518 460046 408574 460102
rect 408642 460046 408698 460102
rect 408518 459922 408574 459978
rect 408642 459922 408698 459978
rect 439238 460294 439294 460350
rect 439362 460294 439418 460350
rect 439238 460170 439294 460226
rect 439362 460170 439418 460226
rect 439238 460046 439294 460102
rect 439362 460046 439418 460102
rect 439238 459922 439294 459978
rect 439362 459922 439418 459978
rect 469958 460294 470014 460350
rect 470082 460294 470138 460350
rect 469958 460170 470014 460226
rect 470082 460170 470138 460226
rect 469958 460046 470014 460102
rect 470082 460046 470138 460102
rect 469958 459922 470014 459978
rect 470082 459922 470138 459978
rect 500678 460294 500734 460350
rect 500802 460294 500858 460350
rect 500678 460170 500734 460226
rect 500802 460170 500858 460226
rect 500678 460046 500734 460102
rect 500802 460046 500858 460102
rect 500678 459922 500734 459978
rect 500802 459922 500858 459978
rect 24518 454294 24574 454350
rect 24642 454294 24698 454350
rect 24518 454170 24574 454226
rect 24642 454170 24698 454226
rect 24518 454046 24574 454102
rect 24642 454046 24698 454102
rect 24518 453922 24574 453978
rect 24642 453922 24698 453978
rect 55238 454294 55294 454350
rect 55362 454294 55418 454350
rect 55238 454170 55294 454226
rect 55362 454170 55418 454226
rect 55238 454046 55294 454102
rect 55362 454046 55418 454102
rect 55238 453922 55294 453978
rect 55362 453922 55418 453978
rect 85958 454294 86014 454350
rect 86082 454294 86138 454350
rect 85958 454170 86014 454226
rect 86082 454170 86138 454226
rect 85958 454046 86014 454102
rect 86082 454046 86138 454102
rect 85958 453922 86014 453978
rect 86082 453922 86138 453978
rect 116678 454294 116734 454350
rect 116802 454294 116858 454350
rect 116678 454170 116734 454226
rect 116802 454170 116858 454226
rect 116678 454046 116734 454102
rect 116802 454046 116858 454102
rect 116678 453922 116734 453978
rect 116802 453922 116858 453978
rect 147398 454294 147454 454350
rect 147522 454294 147578 454350
rect 147398 454170 147454 454226
rect 147522 454170 147578 454226
rect 147398 454046 147454 454102
rect 147522 454046 147578 454102
rect 147398 453922 147454 453978
rect 147522 453922 147578 453978
rect 178118 454294 178174 454350
rect 178242 454294 178298 454350
rect 178118 454170 178174 454226
rect 178242 454170 178298 454226
rect 178118 454046 178174 454102
rect 178242 454046 178298 454102
rect 178118 453922 178174 453978
rect 178242 453922 178298 453978
rect 208838 454294 208894 454350
rect 208962 454294 209018 454350
rect 208838 454170 208894 454226
rect 208962 454170 209018 454226
rect 208838 454046 208894 454102
rect 208962 454046 209018 454102
rect 208838 453922 208894 453978
rect 208962 453922 209018 453978
rect 239558 454294 239614 454350
rect 239682 454294 239738 454350
rect 239558 454170 239614 454226
rect 239682 454170 239738 454226
rect 239558 454046 239614 454102
rect 239682 454046 239738 454102
rect 239558 453922 239614 453978
rect 239682 453922 239738 453978
rect 270278 454294 270334 454350
rect 270402 454294 270458 454350
rect 270278 454170 270334 454226
rect 270402 454170 270458 454226
rect 270278 454046 270334 454102
rect 270402 454046 270458 454102
rect 270278 453922 270334 453978
rect 270402 453922 270458 453978
rect 300998 454294 301054 454350
rect 301122 454294 301178 454350
rect 300998 454170 301054 454226
rect 301122 454170 301178 454226
rect 300998 454046 301054 454102
rect 301122 454046 301178 454102
rect 300998 453922 301054 453978
rect 301122 453922 301178 453978
rect 331718 454294 331774 454350
rect 331842 454294 331898 454350
rect 331718 454170 331774 454226
rect 331842 454170 331898 454226
rect 331718 454046 331774 454102
rect 331842 454046 331898 454102
rect 331718 453922 331774 453978
rect 331842 453922 331898 453978
rect 362438 454294 362494 454350
rect 362562 454294 362618 454350
rect 362438 454170 362494 454226
rect 362562 454170 362618 454226
rect 362438 454046 362494 454102
rect 362562 454046 362618 454102
rect 362438 453922 362494 453978
rect 362562 453922 362618 453978
rect 393158 454294 393214 454350
rect 393282 454294 393338 454350
rect 393158 454170 393214 454226
rect 393282 454170 393338 454226
rect 393158 454046 393214 454102
rect 393282 454046 393338 454102
rect 393158 453922 393214 453978
rect 393282 453922 393338 453978
rect 423878 454294 423934 454350
rect 424002 454294 424058 454350
rect 423878 454170 423934 454226
rect 424002 454170 424058 454226
rect 423878 454046 423934 454102
rect 424002 454046 424058 454102
rect 423878 453922 423934 453978
rect 424002 453922 424058 453978
rect 454598 454294 454654 454350
rect 454722 454294 454778 454350
rect 454598 454170 454654 454226
rect 454722 454170 454778 454226
rect 454598 454046 454654 454102
rect 454722 454046 454778 454102
rect 454598 453922 454654 453978
rect 454722 453922 454778 453978
rect 485318 454294 485374 454350
rect 485442 454294 485498 454350
rect 485318 454170 485374 454226
rect 485442 454170 485498 454226
rect 485318 454046 485374 454102
rect 485442 454046 485498 454102
rect 485318 453922 485374 453978
rect 485442 453922 485498 453978
rect 516038 454294 516094 454350
rect 516162 454294 516218 454350
rect 516038 454170 516094 454226
rect 516162 454170 516218 454226
rect 516038 454046 516094 454102
rect 516162 454046 516218 454102
rect 516038 453922 516094 453978
rect 516162 453922 516218 453978
rect 525250 454294 525306 454350
rect 525374 454294 525430 454350
rect 525498 454294 525554 454350
rect 525622 454294 525678 454350
rect 525250 454170 525306 454226
rect 525374 454170 525430 454226
rect 525498 454170 525554 454226
rect 525622 454170 525678 454226
rect 525250 454046 525306 454102
rect 525374 454046 525430 454102
rect 525498 454046 525554 454102
rect 525622 454046 525678 454102
rect 525250 453922 525306 453978
rect 525374 453922 525430 453978
rect 525498 453922 525554 453978
rect 525622 453922 525678 453978
rect 6970 442294 7026 442350
rect 7094 442294 7150 442350
rect 7218 442294 7274 442350
rect 7342 442294 7398 442350
rect 6970 442170 7026 442226
rect 7094 442170 7150 442226
rect 7218 442170 7274 442226
rect 7342 442170 7398 442226
rect 6970 442046 7026 442102
rect 7094 442046 7150 442102
rect 7218 442046 7274 442102
rect 7342 442046 7398 442102
rect 6970 441922 7026 441978
rect 7094 441922 7150 441978
rect 7218 441922 7274 441978
rect 7342 441922 7398 441978
rect 39878 442294 39934 442350
rect 40002 442294 40058 442350
rect 39878 442170 39934 442226
rect 40002 442170 40058 442226
rect 39878 442046 39934 442102
rect 40002 442046 40058 442102
rect 39878 441922 39934 441978
rect 40002 441922 40058 441978
rect 70598 442294 70654 442350
rect 70722 442294 70778 442350
rect 70598 442170 70654 442226
rect 70722 442170 70778 442226
rect 70598 442046 70654 442102
rect 70722 442046 70778 442102
rect 70598 441922 70654 441978
rect 70722 441922 70778 441978
rect 101318 442294 101374 442350
rect 101442 442294 101498 442350
rect 101318 442170 101374 442226
rect 101442 442170 101498 442226
rect 101318 442046 101374 442102
rect 101442 442046 101498 442102
rect 101318 441922 101374 441978
rect 101442 441922 101498 441978
rect 132038 442294 132094 442350
rect 132162 442294 132218 442350
rect 132038 442170 132094 442226
rect 132162 442170 132218 442226
rect 132038 442046 132094 442102
rect 132162 442046 132218 442102
rect 132038 441922 132094 441978
rect 132162 441922 132218 441978
rect 162758 442294 162814 442350
rect 162882 442294 162938 442350
rect 162758 442170 162814 442226
rect 162882 442170 162938 442226
rect 162758 442046 162814 442102
rect 162882 442046 162938 442102
rect 162758 441922 162814 441978
rect 162882 441922 162938 441978
rect 193478 442294 193534 442350
rect 193602 442294 193658 442350
rect 193478 442170 193534 442226
rect 193602 442170 193658 442226
rect 193478 442046 193534 442102
rect 193602 442046 193658 442102
rect 193478 441922 193534 441978
rect 193602 441922 193658 441978
rect 224198 442294 224254 442350
rect 224322 442294 224378 442350
rect 224198 442170 224254 442226
rect 224322 442170 224378 442226
rect 224198 442046 224254 442102
rect 224322 442046 224378 442102
rect 224198 441922 224254 441978
rect 224322 441922 224378 441978
rect 254918 442294 254974 442350
rect 255042 442294 255098 442350
rect 254918 442170 254974 442226
rect 255042 442170 255098 442226
rect 254918 442046 254974 442102
rect 255042 442046 255098 442102
rect 254918 441922 254974 441978
rect 255042 441922 255098 441978
rect 285638 442294 285694 442350
rect 285762 442294 285818 442350
rect 285638 442170 285694 442226
rect 285762 442170 285818 442226
rect 285638 442046 285694 442102
rect 285762 442046 285818 442102
rect 285638 441922 285694 441978
rect 285762 441922 285818 441978
rect 316358 442294 316414 442350
rect 316482 442294 316538 442350
rect 316358 442170 316414 442226
rect 316482 442170 316538 442226
rect 316358 442046 316414 442102
rect 316482 442046 316538 442102
rect 316358 441922 316414 441978
rect 316482 441922 316538 441978
rect 347078 442294 347134 442350
rect 347202 442294 347258 442350
rect 347078 442170 347134 442226
rect 347202 442170 347258 442226
rect 347078 442046 347134 442102
rect 347202 442046 347258 442102
rect 347078 441922 347134 441978
rect 347202 441922 347258 441978
rect 377798 442294 377854 442350
rect 377922 442294 377978 442350
rect 377798 442170 377854 442226
rect 377922 442170 377978 442226
rect 377798 442046 377854 442102
rect 377922 442046 377978 442102
rect 377798 441922 377854 441978
rect 377922 441922 377978 441978
rect 408518 442294 408574 442350
rect 408642 442294 408698 442350
rect 408518 442170 408574 442226
rect 408642 442170 408698 442226
rect 408518 442046 408574 442102
rect 408642 442046 408698 442102
rect 408518 441922 408574 441978
rect 408642 441922 408698 441978
rect 439238 442294 439294 442350
rect 439362 442294 439418 442350
rect 439238 442170 439294 442226
rect 439362 442170 439418 442226
rect 439238 442046 439294 442102
rect 439362 442046 439418 442102
rect 439238 441922 439294 441978
rect 439362 441922 439418 441978
rect 469958 442294 470014 442350
rect 470082 442294 470138 442350
rect 469958 442170 470014 442226
rect 470082 442170 470138 442226
rect 469958 442046 470014 442102
rect 470082 442046 470138 442102
rect 469958 441922 470014 441978
rect 470082 441922 470138 441978
rect 500678 442294 500734 442350
rect 500802 442294 500858 442350
rect 500678 442170 500734 442226
rect 500802 442170 500858 442226
rect 500678 442046 500734 442102
rect 500802 442046 500858 442102
rect 500678 441922 500734 441978
rect 500802 441922 500858 441978
rect 24518 436294 24574 436350
rect 24642 436294 24698 436350
rect 24518 436170 24574 436226
rect 24642 436170 24698 436226
rect 24518 436046 24574 436102
rect 24642 436046 24698 436102
rect 24518 435922 24574 435978
rect 24642 435922 24698 435978
rect 55238 436294 55294 436350
rect 55362 436294 55418 436350
rect 55238 436170 55294 436226
rect 55362 436170 55418 436226
rect 55238 436046 55294 436102
rect 55362 436046 55418 436102
rect 55238 435922 55294 435978
rect 55362 435922 55418 435978
rect 85958 436294 86014 436350
rect 86082 436294 86138 436350
rect 85958 436170 86014 436226
rect 86082 436170 86138 436226
rect 85958 436046 86014 436102
rect 86082 436046 86138 436102
rect 85958 435922 86014 435978
rect 86082 435922 86138 435978
rect 116678 436294 116734 436350
rect 116802 436294 116858 436350
rect 116678 436170 116734 436226
rect 116802 436170 116858 436226
rect 116678 436046 116734 436102
rect 116802 436046 116858 436102
rect 116678 435922 116734 435978
rect 116802 435922 116858 435978
rect 147398 436294 147454 436350
rect 147522 436294 147578 436350
rect 147398 436170 147454 436226
rect 147522 436170 147578 436226
rect 147398 436046 147454 436102
rect 147522 436046 147578 436102
rect 147398 435922 147454 435978
rect 147522 435922 147578 435978
rect 178118 436294 178174 436350
rect 178242 436294 178298 436350
rect 178118 436170 178174 436226
rect 178242 436170 178298 436226
rect 178118 436046 178174 436102
rect 178242 436046 178298 436102
rect 178118 435922 178174 435978
rect 178242 435922 178298 435978
rect 208838 436294 208894 436350
rect 208962 436294 209018 436350
rect 208838 436170 208894 436226
rect 208962 436170 209018 436226
rect 208838 436046 208894 436102
rect 208962 436046 209018 436102
rect 208838 435922 208894 435978
rect 208962 435922 209018 435978
rect 239558 436294 239614 436350
rect 239682 436294 239738 436350
rect 239558 436170 239614 436226
rect 239682 436170 239738 436226
rect 239558 436046 239614 436102
rect 239682 436046 239738 436102
rect 239558 435922 239614 435978
rect 239682 435922 239738 435978
rect 270278 436294 270334 436350
rect 270402 436294 270458 436350
rect 270278 436170 270334 436226
rect 270402 436170 270458 436226
rect 270278 436046 270334 436102
rect 270402 436046 270458 436102
rect 270278 435922 270334 435978
rect 270402 435922 270458 435978
rect 300998 436294 301054 436350
rect 301122 436294 301178 436350
rect 300998 436170 301054 436226
rect 301122 436170 301178 436226
rect 300998 436046 301054 436102
rect 301122 436046 301178 436102
rect 300998 435922 301054 435978
rect 301122 435922 301178 435978
rect 331718 436294 331774 436350
rect 331842 436294 331898 436350
rect 331718 436170 331774 436226
rect 331842 436170 331898 436226
rect 331718 436046 331774 436102
rect 331842 436046 331898 436102
rect 331718 435922 331774 435978
rect 331842 435922 331898 435978
rect 362438 436294 362494 436350
rect 362562 436294 362618 436350
rect 362438 436170 362494 436226
rect 362562 436170 362618 436226
rect 362438 436046 362494 436102
rect 362562 436046 362618 436102
rect 362438 435922 362494 435978
rect 362562 435922 362618 435978
rect 393158 436294 393214 436350
rect 393282 436294 393338 436350
rect 393158 436170 393214 436226
rect 393282 436170 393338 436226
rect 393158 436046 393214 436102
rect 393282 436046 393338 436102
rect 393158 435922 393214 435978
rect 393282 435922 393338 435978
rect 423878 436294 423934 436350
rect 424002 436294 424058 436350
rect 423878 436170 423934 436226
rect 424002 436170 424058 436226
rect 423878 436046 423934 436102
rect 424002 436046 424058 436102
rect 423878 435922 423934 435978
rect 424002 435922 424058 435978
rect 454598 436294 454654 436350
rect 454722 436294 454778 436350
rect 454598 436170 454654 436226
rect 454722 436170 454778 436226
rect 454598 436046 454654 436102
rect 454722 436046 454778 436102
rect 454598 435922 454654 435978
rect 454722 435922 454778 435978
rect 485318 436294 485374 436350
rect 485442 436294 485498 436350
rect 485318 436170 485374 436226
rect 485442 436170 485498 436226
rect 485318 436046 485374 436102
rect 485442 436046 485498 436102
rect 485318 435922 485374 435978
rect 485442 435922 485498 435978
rect 516038 436294 516094 436350
rect 516162 436294 516218 436350
rect 516038 436170 516094 436226
rect 516162 436170 516218 436226
rect 516038 436046 516094 436102
rect 516162 436046 516218 436102
rect 516038 435922 516094 435978
rect 516162 435922 516218 435978
rect 525250 436294 525306 436350
rect 525374 436294 525430 436350
rect 525498 436294 525554 436350
rect 525622 436294 525678 436350
rect 525250 436170 525306 436226
rect 525374 436170 525430 436226
rect 525498 436170 525554 436226
rect 525622 436170 525678 436226
rect 525250 436046 525306 436102
rect 525374 436046 525430 436102
rect 525498 436046 525554 436102
rect 525622 436046 525678 436102
rect 525250 435922 525306 435978
rect 525374 435922 525430 435978
rect 525498 435922 525554 435978
rect 525622 435922 525678 435978
rect 6970 424294 7026 424350
rect 7094 424294 7150 424350
rect 7218 424294 7274 424350
rect 7342 424294 7398 424350
rect 6970 424170 7026 424226
rect 7094 424170 7150 424226
rect 7218 424170 7274 424226
rect 7342 424170 7398 424226
rect 6970 424046 7026 424102
rect 7094 424046 7150 424102
rect 7218 424046 7274 424102
rect 7342 424046 7398 424102
rect 6970 423922 7026 423978
rect 7094 423922 7150 423978
rect 7218 423922 7274 423978
rect 7342 423922 7398 423978
rect 39878 424294 39934 424350
rect 40002 424294 40058 424350
rect 39878 424170 39934 424226
rect 40002 424170 40058 424226
rect 39878 424046 39934 424102
rect 40002 424046 40058 424102
rect 39878 423922 39934 423978
rect 40002 423922 40058 423978
rect 70598 424294 70654 424350
rect 70722 424294 70778 424350
rect 70598 424170 70654 424226
rect 70722 424170 70778 424226
rect 70598 424046 70654 424102
rect 70722 424046 70778 424102
rect 70598 423922 70654 423978
rect 70722 423922 70778 423978
rect 101318 424294 101374 424350
rect 101442 424294 101498 424350
rect 101318 424170 101374 424226
rect 101442 424170 101498 424226
rect 101318 424046 101374 424102
rect 101442 424046 101498 424102
rect 101318 423922 101374 423978
rect 101442 423922 101498 423978
rect 132038 424294 132094 424350
rect 132162 424294 132218 424350
rect 132038 424170 132094 424226
rect 132162 424170 132218 424226
rect 132038 424046 132094 424102
rect 132162 424046 132218 424102
rect 132038 423922 132094 423978
rect 132162 423922 132218 423978
rect 162758 424294 162814 424350
rect 162882 424294 162938 424350
rect 162758 424170 162814 424226
rect 162882 424170 162938 424226
rect 162758 424046 162814 424102
rect 162882 424046 162938 424102
rect 162758 423922 162814 423978
rect 162882 423922 162938 423978
rect 193478 424294 193534 424350
rect 193602 424294 193658 424350
rect 193478 424170 193534 424226
rect 193602 424170 193658 424226
rect 193478 424046 193534 424102
rect 193602 424046 193658 424102
rect 193478 423922 193534 423978
rect 193602 423922 193658 423978
rect 224198 424294 224254 424350
rect 224322 424294 224378 424350
rect 224198 424170 224254 424226
rect 224322 424170 224378 424226
rect 224198 424046 224254 424102
rect 224322 424046 224378 424102
rect 224198 423922 224254 423978
rect 224322 423922 224378 423978
rect 254918 424294 254974 424350
rect 255042 424294 255098 424350
rect 254918 424170 254974 424226
rect 255042 424170 255098 424226
rect 254918 424046 254974 424102
rect 255042 424046 255098 424102
rect 254918 423922 254974 423978
rect 255042 423922 255098 423978
rect 285638 424294 285694 424350
rect 285762 424294 285818 424350
rect 285638 424170 285694 424226
rect 285762 424170 285818 424226
rect 285638 424046 285694 424102
rect 285762 424046 285818 424102
rect 285638 423922 285694 423978
rect 285762 423922 285818 423978
rect 316358 424294 316414 424350
rect 316482 424294 316538 424350
rect 316358 424170 316414 424226
rect 316482 424170 316538 424226
rect 316358 424046 316414 424102
rect 316482 424046 316538 424102
rect 316358 423922 316414 423978
rect 316482 423922 316538 423978
rect 347078 424294 347134 424350
rect 347202 424294 347258 424350
rect 347078 424170 347134 424226
rect 347202 424170 347258 424226
rect 347078 424046 347134 424102
rect 347202 424046 347258 424102
rect 347078 423922 347134 423978
rect 347202 423922 347258 423978
rect 377798 424294 377854 424350
rect 377922 424294 377978 424350
rect 377798 424170 377854 424226
rect 377922 424170 377978 424226
rect 377798 424046 377854 424102
rect 377922 424046 377978 424102
rect 377798 423922 377854 423978
rect 377922 423922 377978 423978
rect 408518 424294 408574 424350
rect 408642 424294 408698 424350
rect 408518 424170 408574 424226
rect 408642 424170 408698 424226
rect 408518 424046 408574 424102
rect 408642 424046 408698 424102
rect 408518 423922 408574 423978
rect 408642 423922 408698 423978
rect 439238 424294 439294 424350
rect 439362 424294 439418 424350
rect 439238 424170 439294 424226
rect 439362 424170 439418 424226
rect 439238 424046 439294 424102
rect 439362 424046 439418 424102
rect 439238 423922 439294 423978
rect 439362 423922 439418 423978
rect 469958 424294 470014 424350
rect 470082 424294 470138 424350
rect 469958 424170 470014 424226
rect 470082 424170 470138 424226
rect 469958 424046 470014 424102
rect 470082 424046 470138 424102
rect 469958 423922 470014 423978
rect 470082 423922 470138 423978
rect 500678 424294 500734 424350
rect 500802 424294 500858 424350
rect 500678 424170 500734 424226
rect 500802 424170 500858 424226
rect 500678 424046 500734 424102
rect 500802 424046 500858 424102
rect 500678 423922 500734 423978
rect 500802 423922 500858 423978
rect 24518 418294 24574 418350
rect 24642 418294 24698 418350
rect 24518 418170 24574 418226
rect 24642 418170 24698 418226
rect 24518 418046 24574 418102
rect 24642 418046 24698 418102
rect 24518 417922 24574 417978
rect 24642 417922 24698 417978
rect 55238 418294 55294 418350
rect 55362 418294 55418 418350
rect 55238 418170 55294 418226
rect 55362 418170 55418 418226
rect 55238 418046 55294 418102
rect 55362 418046 55418 418102
rect 55238 417922 55294 417978
rect 55362 417922 55418 417978
rect 85958 418294 86014 418350
rect 86082 418294 86138 418350
rect 85958 418170 86014 418226
rect 86082 418170 86138 418226
rect 85958 418046 86014 418102
rect 86082 418046 86138 418102
rect 85958 417922 86014 417978
rect 86082 417922 86138 417978
rect 116678 418294 116734 418350
rect 116802 418294 116858 418350
rect 116678 418170 116734 418226
rect 116802 418170 116858 418226
rect 116678 418046 116734 418102
rect 116802 418046 116858 418102
rect 116678 417922 116734 417978
rect 116802 417922 116858 417978
rect 147398 418294 147454 418350
rect 147522 418294 147578 418350
rect 147398 418170 147454 418226
rect 147522 418170 147578 418226
rect 147398 418046 147454 418102
rect 147522 418046 147578 418102
rect 147398 417922 147454 417978
rect 147522 417922 147578 417978
rect 178118 418294 178174 418350
rect 178242 418294 178298 418350
rect 178118 418170 178174 418226
rect 178242 418170 178298 418226
rect 178118 418046 178174 418102
rect 178242 418046 178298 418102
rect 178118 417922 178174 417978
rect 178242 417922 178298 417978
rect 208838 418294 208894 418350
rect 208962 418294 209018 418350
rect 208838 418170 208894 418226
rect 208962 418170 209018 418226
rect 208838 418046 208894 418102
rect 208962 418046 209018 418102
rect 208838 417922 208894 417978
rect 208962 417922 209018 417978
rect 239558 418294 239614 418350
rect 239682 418294 239738 418350
rect 239558 418170 239614 418226
rect 239682 418170 239738 418226
rect 239558 418046 239614 418102
rect 239682 418046 239738 418102
rect 239558 417922 239614 417978
rect 239682 417922 239738 417978
rect 270278 418294 270334 418350
rect 270402 418294 270458 418350
rect 270278 418170 270334 418226
rect 270402 418170 270458 418226
rect 270278 418046 270334 418102
rect 270402 418046 270458 418102
rect 270278 417922 270334 417978
rect 270402 417922 270458 417978
rect 300998 418294 301054 418350
rect 301122 418294 301178 418350
rect 300998 418170 301054 418226
rect 301122 418170 301178 418226
rect 300998 418046 301054 418102
rect 301122 418046 301178 418102
rect 300998 417922 301054 417978
rect 301122 417922 301178 417978
rect 331718 418294 331774 418350
rect 331842 418294 331898 418350
rect 331718 418170 331774 418226
rect 331842 418170 331898 418226
rect 331718 418046 331774 418102
rect 331842 418046 331898 418102
rect 331718 417922 331774 417978
rect 331842 417922 331898 417978
rect 362438 418294 362494 418350
rect 362562 418294 362618 418350
rect 362438 418170 362494 418226
rect 362562 418170 362618 418226
rect 362438 418046 362494 418102
rect 362562 418046 362618 418102
rect 362438 417922 362494 417978
rect 362562 417922 362618 417978
rect 393158 418294 393214 418350
rect 393282 418294 393338 418350
rect 393158 418170 393214 418226
rect 393282 418170 393338 418226
rect 393158 418046 393214 418102
rect 393282 418046 393338 418102
rect 393158 417922 393214 417978
rect 393282 417922 393338 417978
rect 423878 418294 423934 418350
rect 424002 418294 424058 418350
rect 423878 418170 423934 418226
rect 424002 418170 424058 418226
rect 423878 418046 423934 418102
rect 424002 418046 424058 418102
rect 423878 417922 423934 417978
rect 424002 417922 424058 417978
rect 454598 418294 454654 418350
rect 454722 418294 454778 418350
rect 454598 418170 454654 418226
rect 454722 418170 454778 418226
rect 454598 418046 454654 418102
rect 454722 418046 454778 418102
rect 454598 417922 454654 417978
rect 454722 417922 454778 417978
rect 485318 418294 485374 418350
rect 485442 418294 485498 418350
rect 485318 418170 485374 418226
rect 485442 418170 485498 418226
rect 485318 418046 485374 418102
rect 485442 418046 485498 418102
rect 485318 417922 485374 417978
rect 485442 417922 485498 417978
rect 516038 418294 516094 418350
rect 516162 418294 516218 418350
rect 516038 418170 516094 418226
rect 516162 418170 516218 418226
rect 516038 418046 516094 418102
rect 516162 418046 516218 418102
rect 516038 417922 516094 417978
rect 516162 417922 516218 417978
rect 525250 418294 525306 418350
rect 525374 418294 525430 418350
rect 525498 418294 525554 418350
rect 525622 418294 525678 418350
rect 525250 418170 525306 418226
rect 525374 418170 525430 418226
rect 525498 418170 525554 418226
rect 525622 418170 525678 418226
rect 525250 418046 525306 418102
rect 525374 418046 525430 418102
rect 525498 418046 525554 418102
rect 525622 418046 525678 418102
rect 525250 417922 525306 417978
rect 525374 417922 525430 417978
rect 525498 417922 525554 417978
rect 525622 417922 525678 417978
rect 6970 406294 7026 406350
rect 7094 406294 7150 406350
rect 7218 406294 7274 406350
rect 7342 406294 7398 406350
rect 6970 406170 7026 406226
rect 7094 406170 7150 406226
rect 7218 406170 7274 406226
rect 7342 406170 7398 406226
rect 6970 406046 7026 406102
rect 7094 406046 7150 406102
rect 7218 406046 7274 406102
rect 7342 406046 7398 406102
rect 6970 405922 7026 405978
rect 7094 405922 7150 405978
rect 7218 405922 7274 405978
rect 7342 405922 7398 405978
rect 39878 406294 39934 406350
rect 40002 406294 40058 406350
rect 39878 406170 39934 406226
rect 40002 406170 40058 406226
rect 39878 406046 39934 406102
rect 40002 406046 40058 406102
rect 39878 405922 39934 405978
rect 40002 405922 40058 405978
rect 70598 406294 70654 406350
rect 70722 406294 70778 406350
rect 70598 406170 70654 406226
rect 70722 406170 70778 406226
rect 70598 406046 70654 406102
rect 70722 406046 70778 406102
rect 70598 405922 70654 405978
rect 70722 405922 70778 405978
rect 101318 406294 101374 406350
rect 101442 406294 101498 406350
rect 101318 406170 101374 406226
rect 101442 406170 101498 406226
rect 101318 406046 101374 406102
rect 101442 406046 101498 406102
rect 101318 405922 101374 405978
rect 101442 405922 101498 405978
rect 132038 406294 132094 406350
rect 132162 406294 132218 406350
rect 132038 406170 132094 406226
rect 132162 406170 132218 406226
rect 132038 406046 132094 406102
rect 132162 406046 132218 406102
rect 132038 405922 132094 405978
rect 132162 405922 132218 405978
rect 162758 406294 162814 406350
rect 162882 406294 162938 406350
rect 162758 406170 162814 406226
rect 162882 406170 162938 406226
rect 162758 406046 162814 406102
rect 162882 406046 162938 406102
rect 162758 405922 162814 405978
rect 162882 405922 162938 405978
rect 193478 406294 193534 406350
rect 193602 406294 193658 406350
rect 193478 406170 193534 406226
rect 193602 406170 193658 406226
rect 193478 406046 193534 406102
rect 193602 406046 193658 406102
rect 193478 405922 193534 405978
rect 193602 405922 193658 405978
rect 224198 406294 224254 406350
rect 224322 406294 224378 406350
rect 224198 406170 224254 406226
rect 224322 406170 224378 406226
rect 224198 406046 224254 406102
rect 224322 406046 224378 406102
rect 224198 405922 224254 405978
rect 224322 405922 224378 405978
rect 254918 406294 254974 406350
rect 255042 406294 255098 406350
rect 254918 406170 254974 406226
rect 255042 406170 255098 406226
rect 254918 406046 254974 406102
rect 255042 406046 255098 406102
rect 254918 405922 254974 405978
rect 255042 405922 255098 405978
rect 285638 406294 285694 406350
rect 285762 406294 285818 406350
rect 285638 406170 285694 406226
rect 285762 406170 285818 406226
rect 285638 406046 285694 406102
rect 285762 406046 285818 406102
rect 285638 405922 285694 405978
rect 285762 405922 285818 405978
rect 316358 406294 316414 406350
rect 316482 406294 316538 406350
rect 316358 406170 316414 406226
rect 316482 406170 316538 406226
rect 316358 406046 316414 406102
rect 316482 406046 316538 406102
rect 316358 405922 316414 405978
rect 316482 405922 316538 405978
rect 347078 406294 347134 406350
rect 347202 406294 347258 406350
rect 347078 406170 347134 406226
rect 347202 406170 347258 406226
rect 347078 406046 347134 406102
rect 347202 406046 347258 406102
rect 347078 405922 347134 405978
rect 347202 405922 347258 405978
rect 377798 406294 377854 406350
rect 377922 406294 377978 406350
rect 377798 406170 377854 406226
rect 377922 406170 377978 406226
rect 377798 406046 377854 406102
rect 377922 406046 377978 406102
rect 377798 405922 377854 405978
rect 377922 405922 377978 405978
rect 408518 406294 408574 406350
rect 408642 406294 408698 406350
rect 408518 406170 408574 406226
rect 408642 406170 408698 406226
rect 408518 406046 408574 406102
rect 408642 406046 408698 406102
rect 408518 405922 408574 405978
rect 408642 405922 408698 405978
rect 439238 406294 439294 406350
rect 439362 406294 439418 406350
rect 439238 406170 439294 406226
rect 439362 406170 439418 406226
rect 439238 406046 439294 406102
rect 439362 406046 439418 406102
rect 439238 405922 439294 405978
rect 439362 405922 439418 405978
rect 469958 406294 470014 406350
rect 470082 406294 470138 406350
rect 469958 406170 470014 406226
rect 470082 406170 470138 406226
rect 469958 406046 470014 406102
rect 470082 406046 470138 406102
rect 469958 405922 470014 405978
rect 470082 405922 470138 405978
rect 500678 406294 500734 406350
rect 500802 406294 500858 406350
rect 500678 406170 500734 406226
rect 500802 406170 500858 406226
rect 500678 406046 500734 406102
rect 500802 406046 500858 406102
rect 500678 405922 500734 405978
rect 500802 405922 500858 405978
rect 24518 400294 24574 400350
rect 24642 400294 24698 400350
rect 24518 400170 24574 400226
rect 24642 400170 24698 400226
rect 24518 400046 24574 400102
rect 24642 400046 24698 400102
rect 24518 399922 24574 399978
rect 24642 399922 24698 399978
rect 55238 400294 55294 400350
rect 55362 400294 55418 400350
rect 55238 400170 55294 400226
rect 55362 400170 55418 400226
rect 55238 400046 55294 400102
rect 55362 400046 55418 400102
rect 55238 399922 55294 399978
rect 55362 399922 55418 399978
rect 85958 400294 86014 400350
rect 86082 400294 86138 400350
rect 85958 400170 86014 400226
rect 86082 400170 86138 400226
rect 85958 400046 86014 400102
rect 86082 400046 86138 400102
rect 85958 399922 86014 399978
rect 86082 399922 86138 399978
rect 116678 400294 116734 400350
rect 116802 400294 116858 400350
rect 116678 400170 116734 400226
rect 116802 400170 116858 400226
rect 116678 400046 116734 400102
rect 116802 400046 116858 400102
rect 116678 399922 116734 399978
rect 116802 399922 116858 399978
rect 147398 400294 147454 400350
rect 147522 400294 147578 400350
rect 147398 400170 147454 400226
rect 147522 400170 147578 400226
rect 147398 400046 147454 400102
rect 147522 400046 147578 400102
rect 147398 399922 147454 399978
rect 147522 399922 147578 399978
rect 178118 400294 178174 400350
rect 178242 400294 178298 400350
rect 178118 400170 178174 400226
rect 178242 400170 178298 400226
rect 178118 400046 178174 400102
rect 178242 400046 178298 400102
rect 178118 399922 178174 399978
rect 178242 399922 178298 399978
rect 208838 400294 208894 400350
rect 208962 400294 209018 400350
rect 208838 400170 208894 400226
rect 208962 400170 209018 400226
rect 208838 400046 208894 400102
rect 208962 400046 209018 400102
rect 208838 399922 208894 399978
rect 208962 399922 209018 399978
rect 239558 400294 239614 400350
rect 239682 400294 239738 400350
rect 239558 400170 239614 400226
rect 239682 400170 239738 400226
rect 239558 400046 239614 400102
rect 239682 400046 239738 400102
rect 239558 399922 239614 399978
rect 239682 399922 239738 399978
rect 270278 400294 270334 400350
rect 270402 400294 270458 400350
rect 270278 400170 270334 400226
rect 270402 400170 270458 400226
rect 270278 400046 270334 400102
rect 270402 400046 270458 400102
rect 270278 399922 270334 399978
rect 270402 399922 270458 399978
rect 300998 400294 301054 400350
rect 301122 400294 301178 400350
rect 300998 400170 301054 400226
rect 301122 400170 301178 400226
rect 300998 400046 301054 400102
rect 301122 400046 301178 400102
rect 300998 399922 301054 399978
rect 301122 399922 301178 399978
rect 331718 400294 331774 400350
rect 331842 400294 331898 400350
rect 331718 400170 331774 400226
rect 331842 400170 331898 400226
rect 331718 400046 331774 400102
rect 331842 400046 331898 400102
rect 331718 399922 331774 399978
rect 331842 399922 331898 399978
rect 362438 400294 362494 400350
rect 362562 400294 362618 400350
rect 362438 400170 362494 400226
rect 362562 400170 362618 400226
rect 362438 400046 362494 400102
rect 362562 400046 362618 400102
rect 362438 399922 362494 399978
rect 362562 399922 362618 399978
rect 393158 400294 393214 400350
rect 393282 400294 393338 400350
rect 393158 400170 393214 400226
rect 393282 400170 393338 400226
rect 393158 400046 393214 400102
rect 393282 400046 393338 400102
rect 393158 399922 393214 399978
rect 393282 399922 393338 399978
rect 423878 400294 423934 400350
rect 424002 400294 424058 400350
rect 423878 400170 423934 400226
rect 424002 400170 424058 400226
rect 423878 400046 423934 400102
rect 424002 400046 424058 400102
rect 423878 399922 423934 399978
rect 424002 399922 424058 399978
rect 454598 400294 454654 400350
rect 454722 400294 454778 400350
rect 454598 400170 454654 400226
rect 454722 400170 454778 400226
rect 454598 400046 454654 400102
rect 454722 400046 454778 400102
rect 454598 399922 454654 399978
rect 454722 399922 454778 399978
rect 485318 400294 485374 400350
rect 485442 400294 485498 400350
rect 485318 400170 485374 400226
rect 485442 400170 485498 400226
rect 485318 400046 485374 400102
rect 485442 400046 485498 400102
rect 485318 399922 485374 399978
rect 485442 399922 485498 399978
rect 516038 400294 516094 400350
rect 516162 400294 516218 400350
rect 516038 400170 516094 400226
rect 516162 400170 516218 400226
rect 516038 400046 516094 400102
rect 516162 400046 516218 400102
rect 516038 399922 516094 399978
rect 516162 399922 516218 399978
rect 525250 400294 525306 400350
rect 525374 400294 525430 400350
rect 525498 400294 525554 400350
rect 525622 400294 525678 400350
rect 525250 400170 525306 400226
rect 525374 400170 525430 400226
rect 525498 400170 525554 400226
rect 525622 400170 525678 400226
rect 525250 400046 525306 400102
rect 525374 400046 525430 400102
rect 525498 400046 525554 400102
rect 525622 400046 525678 400102
rect 525250 399922 525306 399978
rect 525374 399922 525430 399978
rect 525498 399922 525554 399978
rect 525622 399922 525678 399978
rect 6970 388294 7026 388350
rect 7094 388294 7150 388350
rect 7218 388294 7274 388350
rect 7342 388294 7398 388350
rect 6970 388170 7026 388226
rect 7094 388170 7150 388226
rect 7218 388170 7274 388226
rect 7342 388170 7398 388226
rect 6970 388046 7026 388102
rect 7094 388046 7150 388102
rect 7218 388046 7274 388102
rect 7342 388046 7398 388102
rect 6970 387922 7026 387978
rect 7094 387922 7150 387978
rect 7218 387922 7274 387978
rect 7342 387922 7398 387978
rect 39878 388294 39934 388350
rect 40002 388294 40058 388350
rect 39878 388170 39934 388226
rect 40002 388170 40058 388226
rect 39878 388046 39934 388102
rect 40002 388046 40058 388102
rect 39878 387922 39934 387978
rect 40002 387922 40058 387978
rect 70598 388294 70654 388350
rect 70722 388294 70778 388350
rect 70598 388170 70654 388226
rect 70722 388170 70778 388226
rect 70598 388046 70654 388102
rect 70722 388046 70778 388102
rect 70598 387922 70654 387978
rect 70722 387922 70778 387978
rect 101318 388294 101374 388350
rect 101442 388294 101498 388350
rect 101318 388170 101374 388226
rect 101442 388170 101498 388226
rect 101318 388046 101374 388102
rect 101442 388046 101498 388102
rect 101318 387922 101374 387978
rect 101442 387922 101498 387978
rect 132038 388294 132094 388350
rect 132162 388294 132218 388350
rect 132038 388170 132094 388226
rect 132162 388170 132218 388226
rect 132038 388046 132094 388102
rect 132162 388046 132218 388102
rect 132038 387922 132094 387978
rect 132162 387922 132218 387978
rect 162758 388294 162814 388350
rect 162882 388294 162938 388350
rect 162758 388170 162814 388226
rect 162882 388170 162938 388226
rect 162758 388046 162814 388102
rect 162882 388046 162938 388102
rect 162758 387922 162814 387978
rect 162882 387922 162938 387978
rect 193478 388294 193534 388350
rect 193602 388294 193658 388350
rect 193478 388170 193534 388226
rect 193602 388170 193658 388226
rect 193478 388046 193534 388102
rect 193602 388046 193658 388102
rect 193478 387922 193534 387978
rect 193602 387922 193658 387978
rect 224198 388294 224254 388350
rect 224322 388294 224378 388350
rect 224198 388170 224254 388226
rect 224322 388170 224378 388226
rect 224198 388046 224254 388102
rect 224322 388046 224378 388102
rect 224198 387922 224254 387978
rect 224322 387922 224378 387978
rect 254918 388294 254974 388350
rect 255042 388294 255098 388350
rect 254918 388170 254974 388226
rect 255042 388170 255098 388226
rect 254918 388046 254974 388102
rect 255042 388046 255098 388102
rect 254918 387922 254974 387978
rect 255042 387922 255098 387978
rect 285638 388294 285694 388350
rect 285762 388294 285818 388350
rect 285638 388170 285694 388226
rect 285762 388170 285818 388226
rect 285638 388046 285694 388102
rect 285762 388046 285818 388102
rect 285638 387922 285694 387978
rect 285762 387922 285818 387978
rect 316358 388294 316414 388350
rect 316482 388294 316538 388350
rect 316358 388170 316414 388226
rect 316482 388170 316538 388226
rect 316358 388046 316414 388102
rect 316482 388046 316538 388102
rect 316358 387922 316414 387978
rect 316482 387922 316538 387978
rect 347078 388294 347134 388350
rect 347202 388294 347258 388350
rect 347078 388170 347134 388226
rect 347202 388170 347258 388226
rect 347078 388046 347134 388102
rect 347202 388046 347258 388102
rect 347078 387922 347134 387978
rect 347202 387922 347258 387978
rect 377798 388294 377854 388350
rect 377922 388294 377978 388350
rect 377798 388170 377854 388226
rect 377922 388170 377978 388226
rect 377798 388046 377854 388102
rect 377922 388046 377978 388102
rect 377798 387922 377854 387978
rect 377922 387922 377978 387978
rect 408518 388294 408574 388350
rect 408642 388294 408698 388350
rect 408518 388170 408574 388226
rect 408642 388170 408698 388226
rect 408518 388046 408574 388102
rect 408642 388046 408698 388102
rect 408518 387922 408574 387978
rect 408642 387922 408698 387978
rect 439238 388294 439294 388350
rect 439362 388294 439418 388350
rect 439238 388170 439294 388226
rect 439362 388170 439418 388226
rect 439238 388046 439294 388102
rect 439362 388046 439418 388102
rect 439238 387922 439294 387978
rect 439362 387922 439418 387978
rect 469958 388294 470014 388350
rect 470082 388294 470138 388350
rect 469958 388170 470014 388226
rect 470082 388170 470138 388226
rect 469958 388046 470014 388102
rect 470082 388046 470138 388102
rect 469958 387922 470014 387978
rect 470082 387922 470138 387978
rect 500678 388294 500734 388350
rect 500802 388294 500858 388350
rect 500678 388170 500734 388226
rect 500802 388170 500858 388226
rect 500678 388046 500734 388102
rect 500802 388046 500858 388102
rect 500678 387922 500734 387978
rect 500802 387922 500858 387978
rect 24518 382294 24574 382350
rect 24642 382294 24698 382350
rect 24518 382170 24574 382226
rect 24642 382170 24698 382226
rect 24518 382046 24574 382102
rect 24642 382046 24698 382102
rect 24518 381922 24574 381978
rect 24642 381922 24698 381978
rect 55238 382294 55294 382350
rect 55362 382294 55418 382350
rect 55238 382170 55294 382226
rect 55362 382170 55418 382226
rect 55238 382046 55294 382102
rect 55362 382046 55418 382102
rect 55238 381922 55294 381978
rect 55362 381922 55418 381978
rect 85958 382294 86014 382350
rect 86082 382294 86138 382350
rect 85958 382170 86014 382226
rect 86082 382170 86138 382226
rect 85958 382046 86014 382102
rect 86082 382046 86138 382102
rect 85958 381922 86014 381978
rect 86082 381922 86138 381978
rect 116678 382294 116734 382350
rect 116802 382294 116858 382350
rect 116678 382170 116734 382226
rect 116802 382170 116858 382226
rect 116678 382046 116734 382102
rect 116802 382046 116858 382102
rect 116678 381922 116734 381978
rect 116802 381922 116858 381978
rect 147398 382294 147454 382350
rect 147522 382294 147578 382350
rect 147398 382170 147454 382226
rect 147522 382170 147578 382226
rect 147398 382046 147454 382102
rect 147522 382046 147578 382102
rect 147398 381922 147454 381978
rect 147522 381922 147578 381978
rect 178118 382294 178174 382350
rect 178242 382294 178298 382350
rect 178118 382170 178174 382226
rect 178242 382170 178298 382226
rect 178118 382046 178174 382102
rect 178242 382046 178298 382102
rect 178118 381922 178174 381978
rect 178242 381922 178298 381978
rect 208838 382294 208894 382350
rect 208962 382294 209018 382350
rect 208838 382170 208894 382226
rect 208962 382170 209018 382226
rect 208838 382046 208894 382102
rect 208962 382046 209018 382102
rect 208838 381922 208894 381978
rect 208962 381922 209018 381978
rect 239558 382294 239614 382350
rect 239682 382294 239738 382350
rect 239558 382170 239614 382226
rect 239682 382170 239738 382226
rect 239558 382046 239614 382102
rect 239682 382046 239738 382102
rect 239558 381922 239614 381978
rect 239682 381922 239738 381978
rect 270278 382294 270334 382350
rect 270402 382294 270458 382350
rect 270278 382170 270334 382226
rect 270402 382170 270458 382226
rect 270278 382046 270334 382102
rect 270402 382046 270458 382102
rect 270278 381922 270334 381978
rect 270402 381922 270458 381978
rect 300998 382294 301054 382350
rect 301122 382294 301178 382350
rect 300998 382170 301054 382226
rect 301122 382170 301178 382226
rect 300998 382046 301054 382102
rect 301122 382046 301178 382102
rect 300998 381922 301054 381978
rect 301122 381922 301178 381978
rect 331718 382294 331774 382350
rect 331842 382294 331898 382350
rect 331718 382170 331774 382226
rect 331842 382170 331898 382226
rect 331718 382046 331774 382102
rect 331842 382046 331898 382102
rect 331718 381922 331774 381978
rect 331842 381922 331898 381978
rect 362438 382294 362494 382350
rect 362562 382294 362618 382350
rect 362438 382170 362494 382226
rect 362562 382170 362618 382226
rect 362438 382046 362494 382102
rect 362562 382046 362618 382102
rect 362438 381922 362494 381978
rect 362562 381922 362618 381978
rect 393158 382294 393214 382350
rect 393282 382294 393338 382350
rect 393158 382170 393214 382226
rect 393282 382170 393338 382226
rect 393158 382046 393214 382102
rect 393282 382046 393338 382102
rect 393158 381922 393214 381978
rect 393282 381922 393338 381978
rect 423878 382294 423934 382350
rect 424002 382294 424058 382350
rect 423878 382170 423934 382226
rect 424002 382170 424058 382226
rect 423878 382046 423934 382102
rect 424002 382046 424058 382102
rect 423878 381922 423934 381978
rect 424002 381922 424058 381978
rect 454598 382294 454654 382350
rect 454722 382294 454778 382350
rect 454598 382170 454654 382226
rect 454722 382170 454778 382226
rect 454598 382046 454654 382102
rect 454722 382046 454778 382102
rect 454598 381922 454654 381978
rect 454722 381922 454778 381978
rect 485318 382294 485374 382350
rect 485442 382294 485498 382350
rect 485318 382170 485374 382226
rect 485442 382170 485498 382226
rect 485318 382046 485374 382102
rect 485442 382046 485498 382102
rect 485318 381922 485374 381978
rect 485442 381922 485498 381978
rect 516038 382294 516094 382350
rect 516162 382294 516218 382350
rect 516038 382170 516094 382226
rect 516162 382170 516218 382226
rect 516038 382046 516094 382102
rect 516162 382046 516218 382102
rect 516038 381922 516094 381978
rect 516162 381922 516218 381978
rect 525250 382294 525306 382350
rect 525374 382294 525430 382350
rect 525498 382294 525554 382350
rect 525622 382294 525678 382350
rect 525250 382170 525306 382226
rect 525374 382170 525430 382226
rect 525498 382170 525554 382226
rect 525622 382170 525678 382226
rect 525250 382046 525306 382102
rect 525374 382046 525430 382102
rect 525498 382046 525554 382102
rect 525622 382046 525678 382102
rect 525250 381922 525306 381978
rect 525374 381922 525430 381978
rect 525498 381922 525554 381978
rect 525622 381922 525678 381978
rect 6970 370294 7026 370350
rect 7094 370294 7150 370350
rect 7218 370294 7274 370350
rect 7342 370294 7398 370350
rect 6970 370170 7026 370226
rect 7094 370170 7150 370226
rect 7218 370170 7274 370226
rect 7342 370170 7398 370226
rect 6970 370046 7026 370102
rect 7094 370046 7150 370102
rect 7218 370046 7274 370102
rect 7342 370046 7398 370102
rect 6970 369922 7026 369978
rect 7094 369922 7150 369978
rect 7218 369922 7274 369978
rect 7342 369922 7398 369978
rect 39878 370294 39934 370350
rect 40002 370294 40058 370350
rect 39878 370170 39934 370226
rect 40002 370170 40058 370226
rect 39878 370046 39934 370102
rect 40002 370046 40058 370102
rect 39878 369922 39934 369978
rect 40002 369922 40058 369978
rect 70598 370294 70654 370350
rect 70722 370294 70778 370350
rect 70598 370170 70654 370226
rect 70722 370170 70778 370226
rect 70598 370046 70654 370102
rect 70722 370046 70778 370102
rect 70598 369922 70654 369978
rect 70722 369922 70778 369978
rect 101318 370294 101374 370350
rect 101442 370294 101498 370350
rect 101318 370170 101374 370226
rect 101442 370170 101498 370226
rect 101318 370046 101374 370102
rect 101442 370046 101498 370102
rect 101318 369922 101374 369978
rect 101442 369922 101498 369978
rect 132038 370294 132094 370350
rect 132162 370294 132218 370350
rect 132038 370170 132094 370226
rect 132162 370170 132218 370226
rect 132038 370046 132094 370102
rect 132162 370046 132218 370102
rect 132038 369922 132094 369978
rect 132162 369922 132218 369978
rect 162758 370294 162814 370350
rect 162882 370294 162938 370350
rect 162758 370170 162814 370226
rect 162882 370170 162938 370226
rect 162758 370046 162814 370102
rect 162882 370046 162938 370102
rect 162758 369922 162814 369978
rect 162882 369922 162938 369978
rect 193478 370294 193534 370350
rect 193602 370294 193658 370350
rect 193478 370170 193534 370226
rect 193602 370170 193658 370226
rect 193478 370046 193534 370102
rect 193602 370046 193658 370102
rect 193478 369922 193534 369978
rect 193602 369922 193658 369978
rect 224198 370294 224254 370350
rect 224322 370294 224378 370350
rect 224198 370170 224254 370226
rect 224322 370170 224378 370226
rect 224198 370046 224254 370102
rect 224322 370046 224378 370102
rect 224198 369922 224254 369978
rect 224322 369922 224378 369978
rect 254918 370294 254974 370350
rect 255042 370294 255098 370350
rect 254918 370170 254974 370226
rect 255042 370170 255098 370226
rect 254918 370046 254974 370102
rect 255042 370046 255098 370102
rect 254918 369922 254974 369978
rect 255042 369922 255098 369978
rect 285638 370294 285694 370350
rect 285762 370294 285818 370350
rect 285638 370170 285694 370226
rect 285762 370170 285818 370226
rect 285638 370046 285694 370102
rect 285762 370046 285818 370102
rect 285638 369922 285694 369978
rect 285762 369922 285818 369978
rect 316358 370294 316414 370350
rect 316482 370294 316538 370350
rect 316358 370170 316414 370226
rect 316482 370170 316538 370226
rect 316358 370046 316414 370102
rect 316482 370046 316538 370102
rect 316358 369922 316414 369978
rect 316482 369922 316538 369978
rect 347078 370294 347134 370350
rect 347202 370294 347258 370350
rect 347078 370170 347134 370226
rect 347202 370170 347258 370226
rect 347078 370046 347134 370102
rect 347202 370046 347258 370102
rect 347078 369922 347134 369978
rect 347202 369922 347258 369978
rect 377798 370294 377854 370350
rect 377922 370294 377978 370350
rect 377798 370170 377854 370226
rect 377922 370170 377978 370226
rect 377798 370046 377854 370102
rect 377922 370046 377978 370102
rect 377798 369922 377854 369978
rect 377922 369922 377978 369978
rect 408518 370294 408574 370350
rect 408642 370294 408698 370350
rect 408518 370170 408574 370226
rect 408642 370170 408698 370226
rect 408518 370046 408574 370102
rect 408642 370046 408698 370102
rect 408518 369922 408574 369978
rect 408642 369922 408698 369978
rect 439238 370294 439294 370350
rect 439362 370294 439418 370350
rect 439238 370170 439294 370226
rect 439362 370170 439418 370226
rect 439238 370046 439294 370102
rect 439362 370046 439418 370102
rect 439238 369922 439294 369978
rect 439362 369922 439418 369978
rect 469958 370294 470014 370350
rect 470082 370294 470138 370350
rect 469958 370170 470014 370226
rect 470082 370170 470138 370226
rect 469958 370046 470014 370102
rect 470082 370046 470138 370102
rect 469958 369922 470014 369978
rect 470082 369922 470138 369978
rect 500678 370294 500734 370350
rect 500802 370294 500858 370350
rect 500678 370170 500734 370226
rect 500802 370170 500858 370226
rect 500678 370046 500734 370102
rect 500802 370046 500858 370102
rect 500678 369922 500734 369978
rect 500802 369922 500858 369978
rect 24518 364294 24574 364350
rect 24642 364294 24698 364350
rect 24518 364170 24574 364226
rect 24642 364170 24698 364226
rect 24518 364046 24574 364102
rect 24642 364046 24698 364102
rect 24518 363922 24574 363978
rect 24642 363922 24698 363978
rect 55238 364294 55294 364350
rect 55362 364294 55418 364350
rect 55238 364170 55294 364226
rect 55362 364170 55418 364226
rect 55238 364046 55294 364102
rect 55362 364046 55418 364102
rect 55238 363922 55294 363978
rect 55362 363922 55418 363978
rect 85958 364294 86014 364350
rect 86082 364294 86138 364350
rect 85958 364170 86014 364226
rect 86082 364170 86138 364226
rect 85958 364046 86014 364102
rect 86082 364046 86138 364102
rect 85958 363922 86014 363978
rect 86082 363922 86138 363978
rect 116678 364294 116734 364350
rect 116802 364294 116858 364350
rect 116678 364170 116734 364226
rect 116802 364170 116858 364226
rect 116678 364046 116734 364102
rect 116802 364046 116858 364102
rect 116678 363922 116734 363978
rect 116802 363922 116858 363978
rect 147398 364294 147454 364350
rect 147522 364294 147578 364350
rect 147398 364170 147454 364226
rect 147522 364170 147578 364226
rect 147398 364046 147454 364102
rect 147522 364046 147578 364102
rect 147398 363922 147454 363978
rect 147522 363922 147578 363978
rect 178118 364294 178174 364350
rect 178242 364294 178298 364350
rect 178118 364170 178174 364226
rect 178242 364170 178298 364226
rect 178118 364046 178174 364102
rect 178242 364046 178298 364102
rect 178118 363922 178174 363978
rect 178242 363922 178298 363978
rect 208838 364294 208894 364350
rect 208962 364294 209018 364350
rect 208838 364170 208894 364226
rect 208962 364170 209018 364226
rect 208838 364046 208894 364102
rect 208962 364046 209018 364102
rect 208838 363922 208894 363978
rect 208962 363922 209018 363978
rect 239558 364294 239614 364350
rect 239682 364294 239738 364350
rect 239558 364170 239614 364226
rect 239682 364170 239738 364226
rect 239558 364046 239614 364102
rect 239682 364046 239738 364102
rect 239558 363922 239614 363978
rect 239682 363922 239738 363978
rect 270278 364294 270334 364350
rect 270402 364294 270458 364350
rect 270278 364170 270334 364226
rect 270402 364170 270458 364226
rect 270278 364046 270334 364102
rect 270402 364046 270458 364102
rect 270278 363922 270334 363978
rect 270402 363922 270458 363978
rect 300998 364294 301054 364350
rect 301122 364294 301178 364350
rect 300998 364170 301054 364226
rect 301122 364170 301178 364226
rect 300998 364046 301054 364102
rect 301122 364046 301178 364102
rect 300998 363922 301054 363978
rect 301122 363922 301178 363978
rect 331718 364294 331774 364350
rect 331842 364294 331898 364350
rect 331718 364170 331774 364226
rect 331842 364170 331898 364226
rect 331718 364046 331774 364102
rect 331842 364046 331898 364102
rect 331718 363922 331774 363978
rect 331842 363922 331898 363978
rect 362438 364294 362494 364350
rect 362562 364294 362618 364350
rect 362438 364170 362494 364226
rect 362562 364170 362618 364226
rect 362438 364046 362494 364102
rect 362562 364046 362618 364102
rect 362438 363922 362494 363978
rect 362562 363922 362618 363978
rect 393158 364294 393214 364350
rect 393282 364294 393338 364350
rect 393158 364170 393214 364226
rect 393282 364170 393338 364226
rect 393158 364046 393214 364102
rect 393282 364046 393338 364102
rect 393158 363922 393214 363978
rect 393282 363922 393338 363978
rect 423878 364294 423934 364350
rect 424002 364294 424058 364350
rect 423878 364170 423934 364226
rect 424002 364170 424058 364226
rect 423878 364046 423934 364102
rect 424002 364046 424058 364102
rect 423878 363922 423934 363978
rect 424002 363922 424058 363978
rect 454598 364294 454654 364350
rect 454722 364294 454778 364350
rect 454598 364170 454654 364226
rect 454722 364170 454778 364226
rect 454598 364046 454654 364102
rect 454722 364046 454778 364102
rect 454598 363922 454654 363978
rect 454722 363922 454778 363978
rect 485318 364294 485374 364350
rect 485442 364294 485498 364350
rect 485318 364170 485374 364226
rect 485442 364170 485498 364226
rect 485318 364046 485374 364102
rect 485442 364046 485498 364102
rect 485318 363922 485374 363978
rect 485442 363922 485498 363978
rect 516038 364294 516094 364350
rect 516162 364294 516218 364350
rect 516038 364170 516094 364226
rect 516162 364170 516218 364226
rect 516038 364046 516094 364102
rect 516162 364046 516218 364102
rect 516038 363922 516094 363978
rect 516162 363922 516218 363978
rect 525250 364294 525306 364350
rect 525374 364294 525430 364350
rect 525498 364294 525554 364350
rect 525622 364294 525678 364350
rect 525250 364170 525306 364226
rect 525374 364170 525430 364226
rect 525498 364170 525554 364226
rect 525622 364170 525678 364226
rect 525250 364046 525306 364102
rect 525374 364046 525430 364102
rect 525498 364046 525554 364102
rect 525622 364046 525678 364102
rect 525250 363922 525306 363978
rect 525374 363922 525430 363978
rect 525498 363922 525554 363978
rect 525622 363922 525678 363978
rect 6970 352294 7026 352350
rect 7094 352294 7150 352350
rect 7218 352294 7274 352350
rect 7342 352294 7398 352350
rect 6970 352170 7026 352226
rect 7094 352170 7150 352226
rect 7218 352170 7274 352226
rect 7342 352170 7398 352226
rect 6970 352046 7026 352102
rect 7094 352046 7150 352102
rect 7218 352046 7274 352102
rect 7342 352046 7398 352102
rect 6970 351922 7026 351978
rect 7094 351922 7150 351978
rect 7218 351922 7274 351978
rect 7342 351922 7398 351978
rect 39878 352294 39934 352350
rect 40002 352294 40058 352350
rect 39878 352170 39934 352226
rect 40002 352170 40058 352226
rect 39878 352046 39934 352102
rect 40002 352046 40058 352102
rect 39878 351922 39934 351978
rect 40002 351922 40058 351978
rect 70598 352294 70654 352350
rect 70722 352294 70778 352350
rect 70598 352170 70654 352226
rect 70722 352170 70778 352226
rect 70598 352046 70654 352102
rect 70722 352046 70778 352102
rect 70598 351922 70654 351978
rect 70722 351922 70778 351978
rect 101318 352294 101374 352350
rect 101442 352294 101498 352350
rect 101318 352170 101374 352226
rect 101442 352170 101498 352226
rect 101318 352046 101374 352102
rect 101442 352046 101498 352102
rect 101318 351922 101374 351978
rect 101442 351922 101498 351978
rect 132038 352294 132094 352350
rect 132162 352294 132218 352350
rect 132038 352170 132094 352226
rect 132162 352170 132218 352226
rect 132038 352046 132094 352102
rect 132162 352046 132218 352102
rect 132038 351922 132094 351978
rect 132162 351922 132218 351978
rect 162758 352294 162814 352350
rect 162882 352294 162938 352350
rect 162758 352170 162814 352226
rect 162882 352170 162938 352226
rect 162758 352046 162814 352102
rect 162882 352046 162938 352102
rect 162758 351922 162814 351978
rect 162882 351922 162938 351978
rect 193478 352294 193534 352350
rect 193602 352294 193658 352350
rect 193478 352170 193534 352226
rect 193602 352170 193658 352226
rect 193478 352046 193534 352102
rect 193602 352046 193658 352102
rect 193478 351922 193534 351978
rect 193602 351922 193658 351978
rect 224198 352294 224254 352350
rect 224322 352294 224378 352350
rect 224198 352170 224254 352226
rect 224322 352170 224378 352226
rect 224198 352046 224254 352102
rect 224322 352046 224378 352102
rect 224198 351922 224254 351978
rect 224322 351922 224378 351978
rect 254918 352294 254974 352350
rect 255042 352294 255098 352350
rect 254918 352170 254974 352226
rect 255042 352170 255098 352226
rect 254918 352046 254974 352102
rect 255042 352046 255098 352102
rect 254918 351922 254974 351978
rect 255042 351922 255098 351978
rect 285638 352294 285694 352350
rect 285762 352294 285818 352350
rect 285638 352170 285694 352226
rect 285762 352170 285818 352226
rect 285638 352046 285694 352102
rect 285762 352046 285818 352102
rect 285638 351922 285694 351978
rect 285762 351922 285818 351978
rect 316358 352294 316414 352350
rect 316482 352294 316538 352350
rect 316358 352170 316414 352226
rect 316482 352170 316538 352226
rect 316358 352046 316414 352102
rect 316482 352046 316538 352102
rect 316358 351922 316414 351978
rect 316482 351922 316538 351978
rect 347078 352294 347134 352350
rect 347202 352294 347258 352350
rect 347078 352170 347134 352226
rect 347202 352170 347258 352226
rect 347078 352046 347134 352102
rect 347202 352046 347258 352102
rect 347078 351922 347134 351978
rect 347202 351922 347258 351978
rect 377798 352294 377854 352350
rect 377922 352294 377978 352350
rect 377798 352170 377854 352226
rect 377922 352170 377978 352226
rect 377798 352046 377854 352102
rect 377922 352046 377978 352102
rect 377798 351922 377854 351978
rect 377922 351922 377978 351978
rect 408518 352294 408574 352350
rect 408642 352294 408698 352350
rect 408518 352170 408574 352226
rect 408642 352170 408698 352226
rect 408518 352046 408574 352102
rect 408642 352046 408698 352102
rect 408518 351922 408574 351978
rect 408642 351922 408698 351978
rect 439238 352294 439294 352350
rect 439362 352294 439418 352350
rect 439238 352170 439294 352226
rect 439362 352170 439418 352226
rect 439238 352046 439294 352102
rect 439362 352046 439418 352102
rect 439238 351922 439294 351978
rect 439362 351922 439418 351978
rect 469958 352294 470014 352350
rect 470082 352294 470138 352350
rect 469958 352170 470014 352226
rect 470082 352170 470138 352226
rect 469958 352046 470014 352102
rect 470082 352046 470138 352102
rect 469958 351922 470014 351978
rect 470082 351922 470138 351978
rect 500678 352294 500734 352350
rect 500802 352294 500858 352350
rect 500678 352170 500734 352226
rect 500802 352170 500858 352226
rect 500678 352046 500734 352102
rect 500802 352046 500858 352102
rect 500678 351922 500734 351978
rect 500802 351922 500858 351978
rect 24518 346294 24574 346350
rect 24642 346294 24698 346350
rect 24518 346170 24574 346226
rect 24642 346170 24698 346226
rect 24518 346046 24574 346102
rect 24642 346046 24698 346102
rect 24518 345922 24574 345978
rect 24642 345922 24698 345978
rect 55238 346294 55294 346350
rect 55362 346294 55418 346350
rect 55238 346170 55294 346226
rect 55362 346170 55418 346226
rect 55238 346046 55294 346102
rect 55362 346046 55418 346102
rect 55238 345922 55294 345978
rect 55362 345922 55418 345978
rect 85958 346294 86014 346350
rect 86082 346294 86138 346350
rect 85958 346170 86014 346226
rect 86082 346170 86138 346226
rect 85958 346046 86014 346102
rect 86082 346046 86138 346102
rect 85958 345922 86014 345978
rect 86082 345922 86138 345978
rect 116678 346294 116734 346350
rect 116802 346294 116858 346350
rect 116678 346170 116734 346226
rect 116802 346170 116858 346226
rect 116678 346046 116734 346102
rect 116802 346046 116858 346102
rect 116678 345922 116734 345978
rect 116802 345922 116858 345978
rect 147398 346294 147454 346350
rect 147522 346294 147578 346350
rect 147398 346170 147454 346226
rect 147522 346170 147578 346226
rect 147398 346046 147454 346102
rect 147522 346046 147578 346102
rect 147398 345922 147454 345978
rect 147522 345922 147578 345978
rect 178118 346294 178174 346350
rect 178242 346294 178298 346350
rect 178118 346170 178174 346226
rect 178242 346170 178298 346226
rect 178118 346046 178174 346102
rect 178242 346046 178298 346102
rect 178118 345922 178174 345978
rect 178242 345922 178298 345978
rect 208838 346294 208894 346350
rect 208962 346294 209018 346350
rect 208838 346170 208894 346226
rect 208962 346170 209018 346226
rect 208838 346046 208894 346102
rect 208962 346046 209018 346102
rect 208838 345922 208894 345978
rect 208962 345922 209018 345978
rect 239558 346294 239614 346350
rect 239682 346294 239738 346350
rect 239558 346170 239614 346226
rect 239682 346170 239738 346226
rect 239558 346046 239614 346102
rect 239682 346046 239738 346102
rect 239558 345922 239614 345978
rect 239682 345922 239738 345978
rect 270278 346294 270334 346350
rect 270402 346294 270458 346350
rect 270278 346170 270334 346226
rect 270402 346170 270458 346226
rect 270278 346046 270334 346102
rect 270402 346046 270458 346102
rect 270278 345922 270334 345978
rect 270402 345922 270458 345978
rect 300998 346294 301054 346350
rect 301122 346294 301178 346350
rect 300998 346170 301054 346226
rect 301122 346170 301178 346226
rect 300998 346046 301054 346102
rect 301122 346046 301178 346102
rect 300998 345922 301054 345978
rect 301122 345922 301178 345978
rect 331718 346294 331774 346350
rect 331842 346294 331898 346350
rect 331718 346170 331774 346226
rect 331842 346170 331898 346226
rect 331718 346046 331774 346102
rect 331842 346046 331898 346102
rect 331718 345922 331774 345978
rect 331842 345922 331898 345978
rect 362438 346294 362494 346350
rect 362562 346294 362618 346350
rect 362438 346170 362494 346226
rect 362562 346170 362618 346226
rect 362438 346046 362494 346102
rect 362562 346046 362618 346102
rect 362438 345922 362494 345978
rect 362562 345922 362618 345978
rect 393158 346294 393214 346350
rect 393282 346294 393338 346350
rect 393158 346170 393214 346226
rect 393282 346170 393338 346226
rect 393158 346046 393214 346102
rect 393282 346046 393338 346102
rect 393158 345922 393214 345978
rect 393282 345922 393338 345978
rect 423878 346294 423934 346350
rect 424002 346294 424058 346350
rect 423878 346170 423934 346226
rect 424002 346170 424058 346226
rect 423878 346046 423934 346102
rect 424002 346046 424058 346102
rect 423878 345922 423934 345978
rect 424002 345922 424058 345978
rect 454598 346294 454654 346350
rect 454722 346294 454778 346350
rect 454598 346170 454654 346226
rect 454722 346170 454778 346226
rect 454598 346046 454654 346102
rect 454722 346046 454778 346102
rect 454598 345922 454654 345978
rect 454722 345922 454778 345978
rect 485318 346294 485374 346350
rect 485442 346294 485498 346350
rect 485318 346170 485374 346226
rect 485442 346170 485498 346226
rect 485318 346046 485374 346102
rect 485442 346046 485498 346102
rect 485318 345922 485374 345978
rect 485442 345922 485498 345978
rect 516038 346294 516094 346350
rect 516162 346294 516218 346350
rect 516038 346170 516094 346226
rect 516162 346170 516218 346226
rect 516038 346046 516094 346102
rect 516162 346046 516218 346102
rect 516038 345922 516094 345978
rect 516162 345922 516218 345978
rect 525250 346294 525306 346350
rect 525374 346294 525430 346350
rect 525498 346294 525554 346350
rect 525622 346294 525678 346350
rect 525250 346170 525306 346226
rect 525374 346170 525430 346226
rect 525498 346170 525554 346226
rect 525622 346170 525678 346226
rect 525250 346046 525306 346102
rect 525374 346046 525430 346102
rect 525498 346046 525554 346102
rect 525622 346046 525678 346102
rect 525250 345922 525306 345978
rect 525374 345922 525430 345978
rect 525498 345922 525554 345978
rect 525622 345922 525678 345978
rect 6970 334294 7026 334350
rect 7094 334294 7150 334350
rect 7218 334294 7274 334350
rect 7342 334294 7398 334350
rect 6970 334170 7026 334226
rect 7094 334170 7150 334226
rect 7218 334170 7274 334226
rect 7342 334170 7398 334226
rect 6970 334046 7026 334102
rect 7094 334046 7150 334102
rect 7218 334046 7274 334102
rect 7342 334046 7398 334102
rect 6970 333922 7026 333978
rect 7094 333922 7150 333978
rect 7218 333922 7274 333978
rect 7342 333922 7398 333978
rect 39878 334294 39934 334350
rect 40002 334294 40058 334350
rect 39878 334170 39934 334226
rect 40002 334170 40058 334226
rect 39878 334046 39934 334102
rect 40002 334046 40058 334102
rect 39878 333922 39934 333978
rect 40002 333922 40058 333978
rect 70598 334294 70654 334350
rect 70722 334294 70778 334350
rect 70598 334170 70654 334226
rect 70722 334170 70778 334226
rect 70598 334046 70654 334102
rect 70722 334046 70778 334102
rect 70598 333922 70654 333978
rect 70722 333922 70778 333978
rect 101318 334294 101374 334350
rect 101442 334294 101498 334350
rect 101318 334170 101374 334226
rect 101442 334170 101498 334226
rect 101318 334046 101374 334102
rect 101442 334046 101498 334102
rect 101318 333922 101374 333978
rect 101442 333922 101498 333978
rect 132038 334294 132094 334350
rect 132162 334294 132218 334350
rect 132038 334170 132094 334226
rect 132162 334170 132218 334226
rect 132038 334046 132094 334102
rect 132162 334046 132218 334102
rect 132038 333922 132094 333978
rect 132162 333922 132218 333978
rect 162758 334294 162814 334350
rect 162882 334294 162938 334350
rect 162758 334170 162814 334226
rect 162882 334170 162938 334226
rect 162758 334046 162814 334102
rect 162882 334046 162938 334102
rect 162758 333922 162814 333978
rect 162882 333922 162938 333978
rect 193478 334294 193534 334350
rect 193602 334294 193658 334350
rect 193478 334170 193534 334226
rect 193602 334170 193658 334226
rect 193478 334046 193534 334102
rect 193602 334046 193658 334102
rect 193478 333922 193534 333978
rect 193602 333922 193658 333978
rect 224198 334294 224254 334350
rect 224322 334294 224378 334350
rect 224198 334170 224254 334226
rect 224322 334170 224378 334226
rect 224198 334046 224254 334102
rect 224322 334046 224378 334102
rect 224198 333922 224254 333978
rect 224322 333922 224378 333978
rect 254918 334294 254974 334350
rect 255042 334294 255098 334350
rect 254918 334170 254974 334226
rect 255042 334170 255098 334226
rect 254918 334046 254974 334102
rect 255042 334046 255098 334102
rect 254918 333922 254974 333978
rect 255042 333922 255098 333978
rect 285638 334294 285694 334350
rect 285762 334294 285818 334350
rect 285638 334170 285694 334226
rect 285762 334170 285818 334226
rect 285638 334046 285694 334102
rect 285762 334046 285818 334102
rect 285638 333922 285694 333978
rect 285762 333922 285818 333978
rect 316358 334294 316414 334350
rect 316482 334294 316538 334350
rect 316358 334170 316414 334226
rect 316482 334170 316538 334226
rect 316358 334046 316414 334102
rect 316482 334046 316538 334102
rect 316358 333922 316414 333978
rect 316482 333922 316538 333978
rect 347078 334294 347134 334350
rect 347202 334294 347258 334350
rect 347078 334170 347134 334226
rect 347202 334170 347258 334226
rect 347078 334046 347134 334102
rect 347202 334046 347258 334102
rect 347078 333922 347134 333978
rect 347202 333922 347258 333978
rect 377798 334294 377854 334350
rect 377922 334294 377978 334350
rect 377798 334170 377854 334226
rect 377922 334170 377978 334226
rect 377798 334046 377854 334102
rect 377922 334046 377978 334102
rect 377798 333922 377854 333978
rect 377922 333922 377978 333978
rect 408518 334294 408574 334350
rect 408642 334294 408698 334350
rect 408518 334170 408574 334226
rect 408642 334170 408698 334226
rect 408518 334046 408574 334102
rect 408642 334046 408698 334102
rect 408518 333922 408574 333978
rect 408642 333922 408698 333978
rect 439238 334294 439294 334350
rect 439362 334294 439418 334350
rect 439238 334170 439294 334226
rect 439362 334170 439418 334226
rect 439238 334046 439294 334102
rect 439362 334046 439418 334102
rect 439238 333922 439294 333978
rect 439362 333922 439418 333978
rect 469958 334294 470014 334350
rect 470082 334294 470138 334350
rect 469958 334170 470014 334226
rect 470082 334170 470138 334226
rect 469958 334046 470014 334102
rect 470082 334046 470138 334102
rect 469958 333922 470014 333978
rect 470082 333922 470138 333978
rect 500678 334294 500734 334350
rect 500802 334294 500858 334350
rect 500678 334170 500734 334226
rect 500802 334170 500858 334226
rect 500678 334046 500734 334102
rect 500802 334046 500858 334102
rect 500678 333922 500734 333978
rect 500802 333922 500858 333978
rect 24518 328294 24574 328350
rect 24642 328294 24698 328350
rect 24518 328170 24574 328226
rect 24642 328170 24698 328226
rect 24518 328046 24574 328102
rect 24642 328046 24698 328102
rect 24518 327922 24574 327978
rect 24642 327922 24698 327978
rect 55238 328294 55294 328350
rect 55362 328294 55418 328350
rect 55238 328170 55294 328226
rect 55362 328170 55418 328226
rect 55238 328046 55294 328102
rect 55362 328046 55418 328102
rect 55238 327922 55294 327978
rect 55362 327922 55418 327978
rect 85958 328294 86014 328350
rect 86082 328294 86138 328350
rect 85958 328170 86014 328226
rect 86082 328170 86138 328226
rect 85958 328046 86014 328102
rect 86082 328046 86138 328102
rect 85958 327922 86014 327978
rect 86082 327922 86138 327978
rect 116678 328294 116734 328350
rect 116802 328294 116858 328350
rect 116678 328170 116734 328226
rect 116802 328170 116858 328226
rect 116678 328046 116734 328102
rect 116802 328046 116858 328102
rect 116678 327922 116734 327978
rect 116802 327922 116858 327978
rect 147398 328294 147454 328350
rect 147522 328294 147578 328350
rect 147398 328170 147454 328226
rect 147522 328170 147578 328226
rect 147398 328046 147454 328102
rect 147522 328046 147578 328102
rect 147398 327922 147454 327978
rect 147522 327922 147578 327978
rect 178118 328294 178174 328350
rect 178242 328294 178298 328350
rect 178118 328170 178174 328226
rect 178242 328170 178298 328226
rect 178118 328046 178174 328102
rect 178242 328046 178298 328102
rect 178118 327922 178174 327978
rect 178242 327922 178298 327978
rect 208838 328294 208894 328350
rect 208962 328294 209018 328350
rect 208838 328170 208894 328226
rect 208962 328170 209018 328226
rect 208838 328046 208894 328102
rect 208962 328046 209018 328102
rect 208838 327922 208894 327978
rect 208962 327922 209018 327978
rect 239558 328294 239614 328350
rect 239682 328294 239738 328350
rect 239558 328170 239614 328226
rect 239682 328170 239738 328226
rect 239558 328046 239614 328102
rect 239682 328046 239738 328102
rect 239558 327922 239614 327978
rect 239682 327922 239738 327978
rect 270278 328294 270334 328350
rect 270402 328294 270458 328350
rect 270278 328170 270334 328226
rect 270402 328170 270458 328226
rect 270278 328046 270334 328102
rect 270402 328046 270458 328102
rect 270278 327922 270334 327978
rect 270402 327922 270458 327978
rect 300998 328294 301054 328350
rect 301122 328294 301178 328350
rect 300998 328170 301054 328226
rect 301122 328170 301178 328226
rect 300998 328046 301054 328102
rect 301122 328046 301178 328102
rect 300998 327922 301054 327978
rect 301122 327922 301178 327978
rect 331718 328294 331774 328350
rect 331842 328294 331898 328350
rect 331718 328170 331774 328226
rect 331842 328170 331898 328226
rect 331718 328046 331774 328102
rect 331842 328046 331898 328102
rect 331718 327922 331774 327978
rect 331842 327922 331898 327978
rect 362438 328294 362494 328350
rect 362562 328294 362618 328350
rect 362438 328170 362494 328226
rect 362562 328170 362618 328226
rect 362438 328046 362494 328102
rect 362562 328046 362618 328102
rect 362438 327922 362494 327978
rect 362562 327922 362618 327978
rect 393158 328294 393214 328350
rect 393282 328294 393338 328350
rect 393158 328170 393214 328226
rect 393282 328170 393338 328226
rect 393158 328046 393214 328102
rect 393282 328046 393338 328102
rect 393158 327922 393214 327978
rect 393282 327922 393338 327978
rect 423878 328294 423934 328350
rect 424002 328294 424058 328350
rect 423878 328170 423934 328226
rect 424002 328170 424058 328226
rect 423878 328046 423934 328102
rect 424002 328046 424058 328102
rect 423878 327922 423934 327978
rect 424002 327922 424058 327978
rect 454598 328294 454654 328350
rect 454722 328294 454778 328350
rect 454598 328170 454654 328226
rect 454722 328170 454778 328226
rect 454598 328046 454654 328102
rect 454722 328046 454778 328102
rect 454598 327922 454654 327978
rect 454722 327922 454778 327978
rect 485318 328294 485374 328350
rect 485442 328294 485498 328350
rect 485318 328170 485374 328226
rect 485442 328170 485498 328226
rect 485318 328046 485374 328102
rect 485442 328046 485498 328102
rect 485318 327922 485374 327978
rect 485442 327922 485498 327978
rect 516038 328294 516094 328350
rect 516162 328294 516218 328350
rect 516038 328170 516094 328226
rect 516162 328170 516218 328226
rect 516038 328046 516094 328102
rect 516162 328046 516218 328102
rect 516038 327922 516094 327978
rect 516162 327922 516218 327978
rect 525250 328294 525306 328350
rect 525374 328294 525430 328350
rect 525498 328294 525554 328350
rect 525622 328294 525678 328350
rect 525250 328170 525306 328226
rect 525374 328170 525430 328226
rect 525498 328170 525554 328226
rect 525622 328170 525678 328226
rect 525250 328046 525306 328102
rect 525374 328046 525430 328102
rect 525498 328046 525554 328102
rect 525622 328046 525678 328102
rect 525250 327922 525306 327978
rect 525374 327922 525430 327978
rect 525498 327922 525554 327978
rect 525622 327922 525678 327978
rect 6970 316294 7026 316350
rect 7094 316294 7150 316350
rect 7218 316294 7274 316350
rect 7342 316294 7398 316350
rect 6970 316170 7026 316226
rect 7094 316170 7150 316226
rect 7218 316170 7274 316226
rect 7342 316170 7398 316226
rect 6970 316046 7026 316102
rect 7094 316046 7150 316102
rect 7218 316046 7274 316102
rect 7342 316046 7398 316102
rect 6970 315922 7026 315978
rect 7094 315922 7150 315978
rect 7218 315922 7274 315978
rect 7342 315922 7398 315978
rect 39878 316294 39934 316350
rect 40002 316294 40058 316350
rect 39878 316170 39934 316226
rect 40002 316170 40058 316226
rect 39878 316046 39934 316102
rect 40002 316046 40058 316102
rect 39878 315922 39934 315978
rect 40002 315922 40058 315978
rect 70598 316294 70654 316350
rect 70722 316294 70778 316350
rect 70598 316170 70654 316226
rect 70722 316170 70778 316226
rect 70598 316046 70654 316102
rect 70722 316046 70778 316102
rect 70598 315922 70654 315978
rect 70722 315922 70778 315978
rect 101318 316294 101374 316350
rect 101442 316294 101498 316350
rect 101318 316170 101374 316226
rect 101442 316170 101498 316226
rect 101318 316046 101374 316102
rect 101442 316046 101498 316102
rect 101318 315922 101374 315978
rect 101442 315922 101498 315978
rect 132038 316294 132094 316350
rect 132162 316294 132218 316350
rect 132038 316170 132094 316226
rect 132162 316170 132218 316226
rect 132038 316046 132094 316102
rect 132162 316046 132218 316102
rect 132038 315922 132094 315978
rect 132162 315922 132218 315978
rect 162758 316294 162814 316350
rect 162882 316294 162938 316350
rect 162758 316170 162814 316226
rect 162882 316170 162938 316226
rect 162758 316046 162814 316102
rect 162882 316046 162938 316102
rect 162758 315922 162814 315978
rect 162882 315922 162938 315978
rect 193478 316294 193534 316350
rect 193602 316294 193658 316350
rect 193478 316170 193534 316226
rect 193602 316170 193658 316226
rect 193478 316046 193534 316102
rect 193602 316046 193658 316102
rect 193478 315922 193534 315978
rect 193602 315922 193658 315978
rect 224198 316294 224254 316350
rect 224322 316294 224378 316350
rect 224198 316170 224254 316226
rect 224322 316170 224378 316226
rect 224198 316046 224254 316102
rect 224322 316046 224378 316102
rect 224198 315922 224254 315978
rect 224322 315922 224378 315978
rect 254918 316294 254974 316350
rect 255042 316294 255098 316350
rect 254918 316170 254974 316226
rect 255042 316170 255098 316226
rect 254918 316046 254974 316102
rect 255042 316046 255098 316102
rect 254918 315922 254974 315978
rect 255042 315922 255098 315978
rect 285638 316294 285694 316350
rect 285762 316294 285818 316350
rect 285638 316170 285694 316226
rect 285762 316170 285818 316226
rect 285638 316046 285694 316102
rect 285762 316046 285818 316102
rect 285638 315922 285694 315978
rect 285762 315922 285818 315978
rect 316358 316294 316414 316350
rect 316482 316294 316538 316350
rect 316358 316170 316414 316226
rect 316482 316170 316538 316226
rect 316358 316046 316414 316102
rect 316482 316046 316538 316102
rect 316358 315922 316414 315978
rect 316482 315922 316538 315978
rect 347078 316294 347134 316350
rect 347202 316294 347258 316350
rect 347078 316170 347134 316226
rect 347202 316170 347258 316226
rect 347078 316046 347134 316102
rect 347202 316046 347258 316102
rect 347078 315922 347134 315978
rect 347202 315922 347258 315978
rect 377798 316294 377854 316350
rect 377922 316294 377978 316350
rect 377798 316170 377854 316226
rect 377922 316170 377978 316226
rect 377798 316046 377854 316102
rect 377922 316046 377978 316102
rect 377798 315922 377854 315978
rect 377922 315922 377978 315978
rect 408518 316294 408574 316350
rect 408642 316294 408698 316350
rect 408518 316170 408574 316226
rect 408642 316170 408698 316226
rect 408518 316046 408574 316102
rect 408642 316046 408698 316102
rect 408518 315922 408574 315978
rect 408642 315922 408698 315978
rect 439238 316294 439294 316350
rect 439362 316294 439418 316350
rect 439238 316170 439294 316226
rect 439362 316170 439418 316226
rect 439238 316046 439294 316102
rect 439362 316046 439418 316102
rect 439238 315922 439294 315978
rect 439362 315922 439418 315978
rect 469958 316294 470014 316350
rect 470082 316294 470138 316350
rect 469958 316170 470014 316226
rect 470082 316170 470138 316226
rect 469958 316046 470014 316102
rect 470082 316046 470138 316102
rect 469958 315922 470014 315978
rect 470082 315922 470138 315978
rect 500678 316294 500734 316350
rect 500802 316294 500858 316350
rect 500678 316170 500734 316226
rect 500802 316170 500858 316226
rect 500678 316046 500734 316102
rect 500802 316046 500858 316102
rect 500678 315922 500734 315978
rect 500802 315922 500858 315978
rect 24518 310294 24574 310350
rect 24642 310294 24698 310350
rect 24518 310170 24574 310226
rect 24642 310170 24698 310226
rect 24518 310046 24574 310102
rect 24642 310046 24698 310102
rect 24518 309922 24574 309978
rect 24642 309922 24698 309978
rect 55238 310294 55294 310350
rect 55362 310294 55418 310350
rect 55238 310170 55294 310226
rect 55362 310170 55418 310226
rect 55238 310046 55294 310102
rect 55362 310046 55418 310102
rect 55238 309922 55294 309978
rect 55362 309922 55418 309978
rect 85958 310294 86014 310350
rect 86082 310294 86138 310350
rect 85958 310170 86014 310226
rect 86082 310170 86138 310226
rect 85958 310046 86014 310102
rect 86082 310046 86138 310102
rect 85958 309922 86014 309978
rect 86082 309922 86138 309978
rect 116678 310294 116734 310350
rect 116802 310294 116858 310350
rect 116678 310170 116734 310226
rect 116802 310170 116858 310226
rect 116678 310046 116734 310102
rect 116802 310046 116858 310102
rect 116678 309922 116734 309978
rect 116802 309922 116858 309978
rect 147398 310294 147454 310350
rect 147522 310294 147578 310350
rect 147398 310170 147454 310226
rect 147522 310170 147578 310226
rect 147398 310046 147454 310102
rect 147522 310046 147578 310102
rect 147398 309922 147454 309978
rect 147522 309922 147578 309978
rect 178118 310294 178174 310350
rect 178242 310294 178298 310350
rect 178118 310170 178174 310226
rect 178242 310170 178298 310226
rect 178118 310046 178174 310102
rect 178242 310046 178298 310102
rect 178118 309922 178174 309978
rect 178242 309922 178298 309978
rect 208838 310294 208894 310350
rect 208962 310294 209018 310350
rect 208838 310170 208894 310226
rect 208962 310170 209018 310226
rect 208838 310046 208894 310102
rect 208962 310046 209018 310102
rect 208838 309922 208894 309978
rect 208962 309922 209018 309978
rect 239558 310294 239614 310350
rect 239682 310294 239738 310350
rect 239558 310170 239614 310226
rect 239682 310170 239738 310226
rect 239558 310046 239614 310102
rect 239682 310046 239738 310102
rect 239558 309922 239614 309978
rect 239682 309922 239738 309978
rect 270278 310294 270334 310350
rect 270402 310294 270458 310350
rect 270278 310170 270334 310226
rect 270402 310170 270458 310226
rect 270278 310046 270334 310102
rect 270402 310046 270458 310102
rect 270278 309922 270334 309978
rect 270402 309922 270458 309978
rect 300998 310294 301054 310350
rect 301122 310294 301178 310350
rect 300998 310170 301054 310226
rect 301122 310170 301178 310226
rect 300998 310046 301054 310102
rect 301122 310046 301178 310102
rect 300998 309922 301054 309978
rect 301122 309922 301178 309978
rect 331718 310294 331774 310350
rect 331842 310294 331898 310350
rect 331718 310170 331774 310226
rect 331842 310170 331898 310226
rect 331718 310046 331774 310102
rect 331842 310046 331898 310102
rect 331718 309922 331774 309978
rect 331842 309922 331898 309978
rect 362438 310294 362494 310350
rect 362562 310294 362618 310350
rect 362438 310170 362494 310226
rect 362562 310170 362618 310226
rect 362438 310046 362494 310102
rect 362562 310046 362618 310102
rect 362438 309922 362494 309978
rect 362562 309922 362618 309978
rect 393158 310294 393214 310350
rect 393282 310294 393338 310350
rect 393158 310170 393214 310226
rect 393282 310170 393338 310226
rect 393158 310046 393214 310102
rect 393282 310046 393338 310102
rect 393158 309922 393214 309978
rect 393282 309922 393338 309978
rect 423878 310294 423934 310350
rect 424002 310294 424058 310350
rect 423878 310170 423934 310226
rect 424002 310170 424058 310226
rect 423878 310046 423934 310102
rect 424002 310046 424058 310102
rect 423878 309922 423934 309978
rect 424002 309922 424058 309978
rect 454598 310294 454654 310350
rect 454722 310294 454778 310350
rect 454598 310170 454654 310226
rect 454722 310170 454778 310226
rect 454598 310046 454654 310102
rect 454722 310046 454778 310102
rect 454598 309922 454654 309978
rect 454722 309922 454778 309978
rect 485318 310294 485374 310350
rect 485442 310294 485498 310350
rect 485318 310170 485374 310226
rect 485442 310170 485498 310226
rect 485318 310046 485374 310102
rect 485442 310046 485498 310102
rect 485318 309922 485374 309978
rect 485442 309922 485498 309978
rect 516038 310294 516094 310350
rect 516162 310294 516218 310350
rect 516038 310170 516094 310226
rect 516162 310170 516218 310226
rect 516038 310046 516094 310102
rect 516162 310046 516218 310102
rect 516038 309922 516094 309978
rect 516162 309922 516218 309978
rect 525250 310294 525306 310350
rect 525374 310294 525430 310350
rect 525498 310294 525554 310350
rect 525622 310294 525678 310350
rect 525250 310170 525306 310226
rect 525374 310170 525430 310226
rect 525498 310170 525554 310226
rect 525622 310170 525678 310226
rect 525250 310046 525306 310102
rect 525374 310046 525430 310102
rect 525498 310046 525554 310102
rect 525622 310046 525678 310102
rect 525250 309922 525306 309978
rect 525374 309922 525430 309978
rect 525498 309922 525554 309978
rect 525622 309922 525678 309978
rect 6970 298294 7026 298350
rect 7094 298294 7150 298350
rect 7218 298294 7274 298350
rect 7342 298294 7398 298350
rect 6970 298170 7026 298226
rect 7094 298170 7150 298226
rect 7218 298170 7274 298226
rect 7342 298170 7398 298226
rect 6970 298046 7026 298102
rect 7094 298046 7150 298102
rect 7218 298046 7274 298102
rect 7342 298046 7398 298102
rect 6970 297922 7026 297978
rect 7094 297922 7150 297978
rect 7218 297922 7274 297978
rect 7342 297922 7398 297978
rect 39878 298294 39934 298350
rect 40002 298294 40058 298350
rect 39878 298170 39934 298226
rect 40002 298170 40058 298226
rect 39878 298046 39934 298102
rect 40002 298046 40058 298102
rect 39878 297922 39934 297978
rect 40002 297922 40058 297978
rect 70598 298294 70654 298350
rect 70722 298294 70778 298350
rect 70598 298170 70654 298226
rect 70722 298170 70778 298226
rect 70598 298046 70654 298102
rect 70722 298046 70778 298102
rect 70598 297922 70654 297978
rect 70722 297922 70778 297978
rect 101318 298294 101374 298350
rect 101442 298294 101498 298350
rect 101318 298170 101374 298226
rect 101442 298170 101498 298226
rect 101318 298046 101374 298102
rect 101442 298046 101498 298102
rect 101318 297922 101374 297978
rect 101442 297922 101498 297978
rect 132038 298294 132094 298350
rect 132162 298294 132218 298350
rect 132038 298170 132094 298226
rect 132162 298170 132218 298226
rect 132038 298046 132094 298102
rect 132162 298046 132218 298102
rect 132038 297922 132094 297978
rect 132162 297922 132218 297978
rect 162758 298294 162814 298350
rect 162882 298294 162938 298350
rect 162758 298170 162814 298226
rect 162882 298170 162938 298226
rect 162758 298046 162814 298102
rect 162882 298046 162938 298102
rect 162758 297922 162814 297978
rect 162882 297922 162938 297978
rect 193478 298294 193534 298350
rect 193602 298294 193658 298350
rect 193478 298170 193534 298226
rect 193602 298170 193658 298226
rect 193478 298046 193534 298102
rect 193602 298046 193658 298102
rect 193478 297922 193534 297978
rect 193602 297922 193658 297978
rect 224198 298294 224254 298350
rect 224322 298294 224378 298350
rect 224198 298170 224254 298226
rect 224322 298170 224378 298226
rect 224198 298046 224254 298102
rect 224322 298046 224378 298102
rect 224198 297922 224254 297978
rect 224322 297922 224378 297978
rect 254918 298294 254974 298350
rect 255042 298294 255098 298350
rect 254918 298170 254974 298226
rect 255042 298170 255098 298226
rect 254918 298046 254974 298102
rect 255042 298046 255098 298102
rect 254918 297922 254974 297978
rect 255042 297922 255098 297978
rect 285638 298294 285694 298350
rect 285762 298294 285818 298350
rect 285638 298170 285694 298226
rect 285762 298170 285818 298226
rect 285638 298046 285694 298102
rect 285762 298046 285818 298102
rect 285638 297922 285694 297978
rect 285762 297922 285818 297978
rect 316358 298294 316414 298350
rect 316482 298294 316538 298350
rect 316358 298170 316414 298226
rect 316482 298170 316538 298226
rect 316358 298046 316414 298102
rect 316482 298046 316538 298102
rect 316358 297922 316414 297978
rect 316482 297922 316538 297978
rect 347078 298294 347134 298350
rect 347202 298294 347258 298350
rect 347078 298170 347134 298226
rect 347202 298170 347258 298226
rect 347078 298046 347134 298102
rect 347202 298046 347258 298102
rect 347078 297922 347134 297978
rect 347202 297922 347258 297978
rect 377798 298294 377854 298350
rect 377922 298294 377978 298350
rect 377798 298170 377854 298226
rect 377922 298170 377978 298226
rect 377798 298046 377854 298102
rect 377922 298046 377978 298102
rect 377798 297922 377854 297978
rect 377922 297922 377978 297978
rect 408518 298294 408574 298350
rect 408642 298294 408698 298350
rect 408518 298170 408574 298226
rect 408642 298170 408698 298226
rect 408518 298046 408574 298102
rect 408642 298046 408698 298102
rect 408518 297922 408574 297978
rect 408642 297922 408698 297978
rect 439238 298294 439294 298350
rect 439362 298294 439418 298350
rect 439238 298170 439294 298226
rect 439362 298170 439418 298226
rect 439238 298046 439294 298102
rect 439362 298046 439418 298102
rect 439238 297922 439294 297978
rect 439362 297922 439418 297978
rect 469958 298294 470014 298350
rect 470082 298294 470138 298350
rect 469958 298170 470014 298226
rect 470082 298170 470138 298226
rect 469958 298046 470014 298102
rect 470082 298046 470138 298102
rect 469958 297922 470014 297978
rect 470082 297922 470138 297978
rect 500678 298294 500734 298350
rect 500802 298294 500858 298350
rect 500678 298170 500734 298226
rect 500802 298170 500858 298226
rect 500678 298046 500734 298102
rect 500802 298046 500858 298102
rect 500678 297922 500734 297978
rect 500802 297922 500858 297978
rect 24518 292294 24574 292350
rect 24642 292294 24698 292350
rect 24518 292170 24574 292226
rect 24642 292170 24698 292226
rect 24518 292046 24574 292102
rect 24642 292046 24698 292102
rect 24518 291922 24574 291978
rect 24642 291922 24698 291978
rect 55238 292294 55294 292350
rect 55362 292294 55418 292350
rect 55238 292170 55294 292226
rect 55362 292170 55418 292226
rect 55238 292046 55294 292102
rect 55362 292046 55418 292102
rect 55238 291922 55294 291978
rect 55362 291922 55418 291978
rect 85958 292294 86014 292350
rect 86082 292294 86138 292350
rect 85958 292170 86014 292226
rect 86082 292170 86138 292226
rect 85958 292046 86014 292102
rect 86082 292046 86138 292102
rect 85958 291922 86014 291978
rect 86082 291922 86138 291978
rect 116678 292294 116734 292350
rect 116802 292294 116858 292350
rect 116678 292170 116734 292226
rect 116802 292170 116858 292226
rect 116678 292046 116734 292102
rect 116802 292046 116858 292102
rect 116678 291922 116734 291978
rect 116802 291922 116858 291978
rect 147398 292294 147454 292350
rect 147522 292294 147578 292350
rect 147398 292170 147454 292226
rect 147522 292170 147578 292226
rect 147398 292046 147454 292102
rect 147522 292046 147578 292102
rect 147398 291922 147454 291978
rect 147522 291922 147578 291978
rect 178118 292294 178174 292350
rect 178242 292294 178298 292350
rect 178118 292170 178174 292226
rect 178242 292170 178298 292226
rect 178118 292046 178174 292102
rect 178242 292046 178298 292102
rect 178118 291922 178174 291978
rect 178242 291922 178298 291978
rect 208838 292294 208894 292350
rect 208962 292294 209018 292350
rect 208838 292170 208894 292226
rect 208962 292170 209018 292226
rect 208838 292046 208894 292102
rect 208962 292046 209018 292102
rect 208838 291922 208894 291978
rect 208962 291922 209018 291978
rect 239558 292294 239614 292350
rect 239682 292294 239738 292350
rect 239558 292170 239614 292226
rect 239682 292170 239738 292226
rect 239558 292046 239614 292102
rect 239682 292046 239738 292102
rect 239558 291922 239614 291978
rect 239682 291922 239738 291978
rect 270278 292294 270334 292350
rect 270402 292294 270458 292350
rect 270278 292170 270334 292226
rect 270402 292170 270458 292226
rect 270278 292046 270334 292102
rect 270402 292046 270458 292102
rect 270278 291922 270334 291978
rect 270402 291922 270458 291978
rect 300998 292294 301054 292350
rect 301122 292294 301178 292350
rect 300998 292170 301054 292226
rect 301122 292170 301178 292226
rect 300998 292046 301054 292102
rect 301122 292046 301178 292102
rect 300998 291922 301054 291978
rect 301122 291922 301178 291978
rect 331718 292294 331774 292350
rect 331842 292294 331898 292350
rect 331718 292170 331774 292226
rect 331842 292170 331898 292226
rect 331718 292046 331774 292102
rect 331842 292046 331898 292102
rect 331718 291922 331774 291978
rect 331842 291922 331898 291978
rect 362438 292294 362494 292350
rect 362562 292294 362618 292350
rect 362438 292170 362494 292226
rect 362562 292170 362618 292226
rect 362438 292046 362494 292102
rect 362562 292046 362618 292102
rect 362438 291922 362494 291978
rect 362562 291922 362618 291978
rect 393158 292294 393214 292350
rect 393282 292294 393338 292350
rect 393158 292170 393214 292226
rect 393282 292170 393338 292226
rect 393158 292046 393214 292102
rect 393282 292046 393338 292102
rect 393158 291922 393214 291978
rect 393282 291922 393338 291978
rect 423878 292294 423934 292350
rect 424002 292294 424058 292350
rect 423878 292170 423934 292226
rect 424002 292170 424058 292226
rect 423878 292046 423934 292102
rect 424002 292046 424058 292102
rect 423878 291922 423934 291978
rect 424002 291922 424058 291978
rect 454598 292294 454654 292350
rect 454722 292294 454778 292350
rect 454598 292170 454654 292226
rect 454722 292170 454778 292226
rect 454598 292046 454654 292102
rect 454722 292046 454778 292102
rect 454598 291922 454654 291978
rect 454722 291922 454778 291978
rect 485318 292294 485374 292350
rect 485442 292294 485498 292350
rect 485318 292170 485374 292226
rect 485442 292170 485498 292226
rect 485318 292046 485374 292102
rect 485442 292046 485498 292102
rect 485318 291922 485374 291978
rect 485442 291922 485498 291978
rect 516038 292294 516094 292350
rect 516162 292294 516218 292350
rect 516038 292170 516094 292226
rect 516162 292170 516218 292226
rect 516038 292046 516094 292102
rect 516162 292046 516218 292102
rect 516038 291922 516094 291978
rect 516162 291922 516218 291978
rect 525250 292294 525306 292350
rect 525374 292294 525430 292350
rect 525498 292294 525554 292350
rect 525622 292294 525678 292350
rect 525250 292170 525306 292226
rect 525374 292170 525430 292226
rect 525498 292170 525554 292226
rect 525622 292170 525678 292226
rect 525250 292046 525306 292102
rect 525374 292046 525430 292102
rect 525498 292046 525554 292102
rect 525622 292046 525678 292102
rect 525250 291922 525306 291978
rect 525374 291922 525430 291978
rect 525498 291922 525554 291978
rect 525622 291922 525678 291978
rect 6970 280294 7026 280350
rect 7094 280294 7150 280350
rect 7218 280294 7274 280350
rect 7342 280294 7398 280350
rect 6970 280170 7026 280226
rect 7094 280170 7150 280226
rect 7218 280170 7274 280226
rect 7342 280170 7398 280226
rect 6970 280046 7026 280102
rect 7094 280046 7150 280102
rect 7218 280046 7274 280102
rect 7342 280046 7398 280102
rect 6970 279922 7026 279978
rect 7094 279922 7150 279978
rect 7218 279922 7274 279978
rect 7342 279922 7398 279978
rect 39878 280294 39934 280350
rect 40002 280294 40058 280350
rect 39878 280170 39934 280226
rect 40002 280170 40058 280226
rect 39878 280046 39934 280102
rect 40002 280046 40058 280102
rect 39878 279922 39934 279978
rect 40002 279922 40058 279978
rect 70598 280294 70654 280350
rect 70722 280294 70778 280350
rect 70598 280170 70654 280226
rect 70722 280170 70778 280226
rect 70598 280046 70654 280102
rect 70722 280046 70778 280102
rect 70598 279922 70654 279978
rect 70722 279922 70778 279978
rect 101318 280294 101374 280350
rect 101442 280294 101498 280350
rect 101318 280170 101374 280226
rect 101442 280170 101498 280226
rect 101318 280046 101374 280102
rect 101442 280046 101498 280102
rect 101318 279922 101374 279978
rect 101442 279922 101498 279978
rect 132038 280294 132094 280350
rect 132162 280294 132218 280350
rect 132038 280170 132094 280226
rect 132162 280170 132218 280226
rect 132038 280046 132094 280102
rect 132162 280046 132218 280102
rect 132038 279922 132094 279978
rect 132162 279922 132218 279978
rect 162758 280294 162814 280350
rect 162882 280294 162938 280350
rect 162758 280170 162814 280226
rect 162882 280170 162938 280226
rect 162758 280046 162814 280102
rect 162882 280046 162938 280102
rect 162758 279922 162814 279978
rect 162882 279922 162938 279978
rect 193478 280294 193534 280350
rect 193602 280294 193658 280350
rect 193478 280170 193534 280226
rect 193602 280170 193658 280226
rect 193478 280046 193534 280102
rect 193602 280046 193658 280102
rect 193478 279922 193534 279978
rect 193602 279922 193658 279978
rect 224198 280294 224254 280350
rect 224322 280294 224378 280350
rect 224198 280170 224254 280226
rect 224322 280170 224378 280226
rect 224198 280046 224254 280102
rect 224322 280046 224378 280102
rect 224198 279922 224254 279978
rect 224322 279922 224378 279978
rect 254918 280294 254974 280350
rect 255042 280294 255098 280350
rect 254918 280170 254974 280226
rect 255042 280170 255098 280226
rect 254918 280046 254974 280102
rect 255042 280046 255098 280102
rect 254918 279922 254974 279978
rect 255042 279922 255098 279978
rect 285638 280294 285694 280350
rect 285762 280294 285818 280350
rect 285638 280170 285694 280226
rect 285762 280170 285818 280226
rect 285638 280046 285694 280102
rect 285762 280046 285818 280102
rect 285638 279922 285694 279978
rect 285762 279922 285818 279978
rect 316358 280294 316414 280350
rect 316482 280294 316538 280350
rect 316358 280170 316414 280226
rect 316482 280170 316538 280226
rect 316358 280046 316414 280102
rect 316482 280046 316538 280102
rect 316358 279922 316414 279978
rect 316482 279922 316538 279978
rect 347078 280294 347134 280350
rect 347202 280294 347258 280350
rect 347078 280170 347134 280226
rect 347202 280170 347258 280226
rect 347078 280046 347134 280102
rect 347202 280046 347258 280102
rect 347078 279922 347134 279978
rect 347202 279922 347258 279978
rect 377798 280294 377854 280350
rect 377922 280294 377978 280350
rect 377798 280170 377854 280226
rect 377922 280170 377978 280226
rect 377798 280046 377854 280102
rect 377922 280046 377978 280102
rect 377798 279922 377854 279978
rect 377922 279922 377978 279978
rect 408518 280294 408574 280350
rect 408642 280294 408698 280350
rect 408518 280170 408574 280226
rect 408642 280170 408698 280226
rect 408518 280046 408574 280102
rect 408642 280046 408698 280102
rect 408518 279922 408574 279978
rect 408642 279922 408698 279978
rect 439238 280294 439294 280350
rect 439362 280294 439418 280350
rect 439238 280170 439294 280226
rect 439362 280170 439418 280226
rect 439238 280046 439294 280102
rect 439362 280046 439418 280102
rect 439238 279922 439294 279978
rect 439362 279922 439418 279978
rect 469958 280294 470014 280350
rect 470082 280294 470138 280350
rect 469958 280170 470014 280226
rect 470082 280170 470138 280226
rect 469958 280046 470014 280102
rect 470082 280046 470138 280102
rect 469958 279922 470014 279978
rect 470082 279922 470138 279978
rect 500678 280294 500734 280350
rect 500802 280294 500858 280350
rect 500678 280170 500734 280226
rect 500802 280170 500858 280226
rect 500678 280046 500734 280102
rect 500802 280046 500858 280102
rect 500678 279922 500734 279978
rect 500802 279922 500858 279978
rect 24518 274294 24574 274350
rect 24642 274294 24698 274350
rect 24518 274170 24574 274226
rect 24642 274170 24698 274226
rect 24518 274046 24574 274102
rect 24642 274046 24698 274102
rect 24518 273922 24574 273978
rect 24642 273922 24698 273978
rect 55238 274294 55294 274350
rect 55362 274294 55418 274350
rect 55238 274170 55294 274226
rect 55362 274170 55418 274226
rect 55238 274046 55294 274102
rect 55362 274046 55418 274102
rect 55238 273922 55294 273978
rect 55362 273922 55418 273978
rect 85958 274294 86014 274350
rect 86082 274294 86138 274350
rect 85958 274170 86014 274226
rect 86082 274170 86138 274226
rect 85958 274046 86014 274102
rect 86082 274046 86138 274102
rect 85958 273922 86014 273978
rect 86082 273922 86138 273978
rect 116678 274294 116734 274350
rect 116802 274294 116858 274350
rect 116678 274170 116734 274226
rect 116802 274170 116858 274226
rect 116678 274046 116734 274102
rect 116802 274046 116858 274102
rect 116678 273922 116734 273978
rect 116802 273922 116858 273978
rect 147398 274294 147454 274350
rect 147522 274294 147578 274350
rect 147398 274170 147454 274226
rect 147522 274170 147578 274226
rect 147398 274046 147454 274102
rect 147522 274046 147578 274102
rect 147398 273922 147454 273978
rect 147522 273922 147578 273978
rect 178118 274294 178174 274350
rect 178242 274294 178298 274350
rect 178118 274170 178174 274226
rect 178242 274170 178298 274226
rect 178118 274046 178174 274102
rect 178242 274046 178298 274102
rect 178118 273922 178174 273978
rect 178242 273922 178298 273978
rect 208838 274294 208894 274350
rect 208962 274294 209018 274350
rect 208838 274170 208894 274226
rect 208962 274170 209018 274226
rect 208838 274046 208894 274102
rect 208962 274046 209018 274102
rect 208838 273922 208894 273978
rect 208962 273922 209018 273978
rect 239558 274294 239614 274350
rect 239682 274294 239738 274350
rect 239558 274170 239614 274226
rect 239682 274170 239738 274226
rect 239558 274046 239614 274102
rect 239682 274046 239738 274102
rect 239558 273922 239614 273978
rect 239682 273922 239738 273978
rect 270278 274294 270334 274350
rect 270402 274294 270458 274350
rect 270278 274170 270334 274226
rect 270402 274170 270458 274226
rect 270278 274046 270334 274102
rect 270402 274046 270458 274102
rect 270278 273922 270334 273978
rect 270402 273922 270458 273978
rect 300998 274294 301054 274350
rect 301122 274294 301178 274350
rect 300998 274170 301054 274226
rect 301122 274170 301178 274226
rect 300998 274046 301054 274102
rect 301122 274046 301178 274102
rect 300998 273922 301054 273978
rect 301122 273922 301178 273978
rect 331718 274294 331774 274350
rect 331842 274294 331898 274350
rect 331718 274170 331774 274226
rect 331842 274170 331898 274226
rect 331718 274046 331774 274102
rect 331842 274046 331898 274102
rect 331718 273922 331774 273978
rect 331842 273922 331898 273978
rect 362438 274294 362494 274350
rect 362562 274294 362618 274350
rect 362438 274170 362494 274226
rect 362562 274170 362618 274226
rect 362438 274046 362494 274102
rect 362562 274046 362618 274102
rect 362438 273922 362494 273978
rect 362562 273922 362618 273978
rect 393158 274294 393214 274350
rect 393282 274294 393338 274350
rect 393158 274170 393214 274226
rect 393282 274170 393338 274226
rect 393158 274046 393214 274102
rect 393282 274046 393338 274102
rect 393158 273922 393214 273978
rect 393282 273922 393338 273978
rect 423878 274294 423934 274350
rect 424002 274294 424058 274350
rect 423878 274170 423934 274226
rect 424002 274170 424058 274226
rect 423878 274046 423934 274102
rect 424002 274046 424058 274102
rect 423878 273922 423934 273978
rect 424002 273922 424058 273978
rect 454598 274294 454654 274350
rect 454722 274294 454778 274350
rect 454598 274170 454654 274226
rect 454722 274170 454778 274226
rect 454598 274046 454654 274102
rect 454722 274046 454778 274102
rect 454598 273922 454654 273978
rect 454722 273922 454778 273978
rect 485318 274294 485374 274350
rect 485442 274294 485498 274350
rect 485318 274170 485374 274226
rect 485442 274170 485498 274226
rect 485318 274046 485374 274102
rect 485442 274046 485498 274102
rect 485318 273922 485374 273978
rect 485442 273922 485498 273978
rect 516038 274294 516094 274350
rect 516162 274294 516218 274350
rect 516038 274170 516094 274226
rect 516162 274170 516218 274226
rect 516038 274046 516094 274102
rect 516162 274046 516218 274102
rect 516038 273922 516094 273978
rect 516162 273922 516218 273978
rect 525250 274294 525306 274350
rect 525374 274294 525430 274350
rect 525498 274294 525554 274350
rect 525622 274294 525678 274350
rect 525250 274170 525306 274226
rect 525374 274170 525430 274226
rect 525498 274170 525554 274226
rect 525622 274170 525678 274226
rect 525250 274046 525306 274102
rect 525374 274046 525430 274102
rect 525498 274046 525554 274102
rect 525622 274046 525678 274102
rect 525250 273922 525306 273978
rect 525374 273922 525430 273978
rect 525498 273922 525554 273978
rect 525622 273922 525678 273978
rect 6970 262294 7026 262350
rect 7094 262294 7150 262350
rect 7218 262294 7274 262350
rect 7342 262294 7398 262350
rect 6970 262170 7026 262226
rect 7094 262170 7150 262226
rect 7218 262170 7274 262226
rect 7342 262170 7398 262226
rect 6970 262046 7026 262102
rect 7094 262046 7150 262102
rect 7218 262046 7274 262102
rect 7342 262046 7398 262102
rect 6970 261922 7026 261978
rect 7094 261922 7150 261978
rect 7218 261922 7274 261978
rect 7342 261922 7398 261978
rect 39878 262294 39934 262350
rect 40002 262294 40058 262350
rect 39878 262170 39934 262226
rect 40002 262170 40058 262226
rect 39878 262046 39934 262102
rect 40002 262046 40058 262102
rect 39878 261922 39934 261978
rect 40002 261922 40058 261978
rect 70598 262294 70654 262350
rect 70722 262294 70778 262350
rect 70598 262170 70654 262226
rect 70722 262170 70778 262226
rect 70598 262046 70654 262102
rect 70722 262046 70778 262102
rect 70598 261922 70654 261978
rect 70722 261922 70778 261978
rect 101318 262294 101374 262350
rect 101442 262294 101498 262350
rect 101318 262170 101374 262226
rect 101442 262170 101498 262226
rect 101318 262046 101374 262102
rect 101442 262046 101498 262102
rect 101318 261922 101374 261978
rect 101442 261922 101498 261978
rect 132038 262294 132094 262350
rect 132162 262294 132218 262350
rect 132038 262170 132094 262226
rect 132162 262170 132218 262226
rect 132038 262046 132094 262102
rect 132162 262046 132218 262102
rect 132038 261922 132094 261978
rect 132162 261922 132218 261978
rect 162758 262294 162814 262350
rect 162882 262294 162938 262350
rect 162758 262170 162814 262226
rect 162882 262170 162938 262226
rect 162758 262046 162814 262102
rect 162882 262046 162938 262102
rect 162758 261922 162814 261978
rect 162882 261922 162938 261978
rect 193478 262294 193534 262350
rect 193602 262294 193658 262350
rect 193478 262170 193534 262226
rect 193602 262170 193658 262226
rect 193478 262046 193534 262102
rect 193602 262046 193658 262102
rect 193478 261922 193534 261978
rect 193602 261922 193658 261978
rect 224198 262294 224254 262350
rect 224322 262294 224378 262350
rect 224198 262170 224254 262226
rect 224322 262170 224378 262226
rect 224198 262046 224254 262102
rect 224322 262046 224378 262102
rect 224198 261922 224254 261978
rect 224322 261922 224378 261978
rect 254918 262294 254974 262350
rect 255042 262294 255098 262350
rect 254918 262170 254974 262226
rect 255042 262170 255098 262226
rect 254918 262046 254974 262102
rect 255042 262046 255098 262102
rect 254918 261922 254974 261978
rect 255042 261922 255098 261978
rect 285638 262294 285694 262350
rect 285762 262294 285818 262350
rect 285638 262170 285694 262226
rect 285762 262170 285818 262226
rect 285638 262046 285694 262102
rect 285762 262046 285818 262102
rect 285638 261922 285694 261978
rect 285762 261922 285818 261978
rect 316358 262294 316414 262350
rect 316482 262294 316538 262350
rect 316358 262170 316414 262226
rect 316482 262170 316538 262226
rect 316358 262046 316414 262102
rect 316482 262046 316538 262102
rect 316358 261922 316414 261978
rect 316482 261922 316538 261978
rect 347078 262294 347134 262350
rect 347202 262294 347258 262350
rect 347078 262170 347134 262226
rect 347202 262170 347258 262226
rect 347078 262046 347134 262102
rect 347202 262046 347258 262102
rect 347078 261922 347134 261978
rect 347202 261922 347258 261978
rect 377798 262294 377854 262350
rect 377922 262294 377978 262350
rect 377798 262170 377854 262226
rect 377922 262170 377978 262226
rect 377798 262046 377854 262102
rect 377922 262046 377978 262102
rect 377798 261922 377854 261978
rect 377922 261922 377978 261978
rect 408518 262294 408574 262350
rect 408642 262294 408698 262350
rect 408518 262170 408574 262226
rect 408642 262170 408698 262226
rect 408518 262046 408574 262102
rect 408642 262046 408698 262102
rect 408518 261922 408574 261978
rect 408642 261922 408698 261978
rect 439238 262294 439294 262350
rect 439362 262294 439418 262350
rect 439238 262170 439294 262226
rect 439362 262170 439418 262226
rect 439238 262046 439294 262102
rect 439362 262046 439418 262102
rect 439238 261922 439294 261978
rect 439362 261922 439418 261978
rect 469958 262294 470014 262350
rect 470082 262294 470138 262350
rect 469958 262170 470014 262226
rect 470082 262170 470138 262226
rect 469958 262046 470014 262102
rect 470082 262046 470138 262102
rect 469958 261922 470014 261978
rect 470082 261922 470138 261978
rect 500678 262294 500734 262350
rect 500802 262294 500858 262350
rect 500678 262170 500734 262226
rect 500802 262170 500858 262226
rect 500678 262046 500734 262102
rect 500802 262046 500858 262102
rect 500678 261922 500734 261978
rect 500802 261922 500858 261978
rect 24518 256294 24574 256350
rect 24642 256294 24698 256350
rect 24518 256170 24574 256226
rect 24642 256170 24698 256226
rect 24518 256046 24574 256102
rect 24642 256046 24698 256102
rect 24518 255922 24574 255978
rect 24642 255922 24698 255978
rect 55238 256294 55294 256350
rect 55362 256294 55418 256350
rect 55238 256170 55294 256226
rect 55362 256170 55418 256226
rect 55238 256046 55294 256102
rect 55362 256046 55418 256102
rect 55238 255922 55294 255978
rect 55362 255922 55418 255978
rect 85958 256294 86014 256350
rect 86082 256294 86138 256350
rect 85958 256170 86014 256226
rect 86082 256170 86138 256226
rect 85958 256046 86014 256102
rect 86082 256046 86138 256102
rect 85958 255922 86014 255978
rect 86082 255922 86138 255978
rect 116678 256294 116734 256350
rect 116802 256294 116858 256350
rect 116678 256170 116734 256226
rect 116802 256170 116858 256226
rect 116678 256046 116734 256102
rect 116802 256046 116858 256102
rect 116678 255922 116734 255978
rect 116802 255922 116858 255978
rect 147398 256294 147454 256350
rect 147522 256294 147578 256350
rect 147398 256170 147454 256226
rect 147522 256170 147578 256226
rect 147398 256046 147454 256102
rect 147522 256046 147578 256102
rect 147398 255922 147454 255978
rect 147522 255922 147578 255978
rect 178118 256294 178174 256350
rect 178242 256294 178298 256350
rect 178118 256170 178174 256226
rect 178242 256170 178298 256226
rect 178118 256046 178174 256102
rect 178242 256046 178298 256102
rect 178118 255922 178174 255978
rect 178242 255922 178298 255978
rect 208838 256294 208894 256350
rect 208962 256294 209018 256350
rect 208838 256170 208894 256226
rect 208962 256170 209018 256226
rect 208838 256046 208894 256102
rect 208962 256046 209018 256102
rect 208838 255922 208894 255978
rect 208962 255922 209018 255978
rect 239558 256294 239614 256350
rect 239682 256294 239738 256350
rect 239558 256170 239614 256226
rect 239682 256170 239738 256226
rect 239558 256046 239614 256102
rect 239682 256046 239738 256102
rect 239558 255922 239614 255978
rect 239682 255922 239738 255978
rect 270278 256294 270334 256350
rect 270402 256294 270458 256350
rect 270278 256170 270334 256226
rect 270402 256170 270458 256226
rect 270278 256046 270334 256102
rect 270402 256046 270458 256102
rect 270278 255922 270334 255978
rect 270402 255922 270458 255978
rect 300998 256294 301054 256350
rect 301122 256294 301178 256350
rect 300998 256170 301054 256226
rect 301122 256170 301178 256226
rect 300998 256046 301054 256102
rect 301122 256046 301178 256102
rect 300998 255922 301054 255978
rect 301122 255922 301178 255978
rect 331718 256294 331774 256350
rect 331842 256294 331898 256350
rect 331718 256170 331774 256226
rect 331842 256170 331898 256226
rect 331718 256046 331774 256102
rect 331842 256046 331898 256102
rect 331718 255922 331774 255978
rect 331842 255922 331898 255978
rect 362438 256294 362494 256350
rect 362562 256294 362618 256350
rect 362438 256170 362494 256226
rect 362562 256170 362618 256226
rect 362438 256046 362494 256102
rect 362562 256046 362618 256102
rect 362438 255922 362494 255978
rect 362562 255922 362618 255978
rect 393158 256294 393214 256350
rect 393282 256294 393338 256350
rect 393158 256170 393214 256226
rect 393282 256170 393338 256226
rect 393158 256046 393214 256102
rect 393282 256046 393338 256102
rect 393158 255922 393214 255978
rect 393282 255922 393338 255978
rect 423878 256294 423934 256350
rect 424002 256294 424058 256350
rect 423878 256170 423934 256226
rect 424002 256170 424058 256226
rect 423878 256046 423934 256102
rect 424002 256046 424058 256102
rect 423878 255922 423934 255978
rect 424002 255922 424058 255978
rect 454598 256294 454654 256350
rect 454722 256294 454778 256350
rect 454598 256170 454654 256226
rect 454722 256170 454778 256226
rect 454598 256046 454654 256102
rect 454722 256046 454778 256102
rect 454598 255922 454654 255978
rect 454722 255922 454778 255978
rect 485318 256294 485374 256350
rect 485442 256294 485498 256350
rect 485318 256170 485374 256226
rect 485442 256170 485498 256226
rect 485318 256046 485374 256102
rect 485442 256046 485498 256102
rect 485318 255922 485374 255978
rect 485442 255922 485498 255978
rect 516038 256294 516094 256350
rect 516162 256294 516218 256350
rect 516038 256170 516094 256226
rect 516162 256170 516218 256226
rect 516038 256046 516094 256102
rect 516162 256046 516218 256102
rect 516038 255922 516094 255978
rect 516162 255922 516218 255978
rect 525250 256294 525306 256350
rect 525374 256294 525430 256350
rect 525498 256294 525554 256350
rect 525622 256294 525678 256350
rect 525250 256170 525306 256226
rect 525374 256170 525430 256226
rect 525498 256170 525554 256226
rect 525622 256170 525678 256226
rect 525250 256046 525306 256102
rect 525374 256046 525430 256102
rect 525498 256046 525554 256102
rect 525622 256046 525678 256102
rect 525250 255922 525306 255978
rect 525374 255922 525430 255978
rect 525498 255922 525554 255978
rect 525622 255922 525678 255978
rect 6970 244294 7026 244350
rect 7094 244294 7150 244350
rect 7218 244294 7274 244350
rect 7342 244294 7398 244350
rect 6970 244170 7026 244226
rect 7094 244170 7150 244226
rect 7218 244170 7274 244226
rect 7342 244170 7398 244226
rect 6970 244046 7026 244102
rect 7094 244046 7150 244102
rect 7218 244046 7274 244102
rect 7342 244046 7398 244102
rect 6970 243922 7026 243978
rect 7094 243922 7150 243978
rect 7218 243922 7274 243978
rect 7342 243922 7398 243978
rect 39878 244294 39934 244350
rect 40002 244294 40058 244350
rect 39878 244170 39934 244226
rect 40002 244170 40058 244226
rect 39878 244046 39934 244102
rect 40002 244046 40058 244102
rect 39878 243922 39934 243978
rect 40002 243922 40058 243978
rect 70598 244294 70654 244350
rect 70722 244294 70778 244350
rect 70598 244170 70654 244226
rect 70722 244170 70778 244226
rect 70598 244046 70654 244102
rect 70722 244046 70778 244102
rect 70598 243922 70654 243978
rect 70722 243922 70778 243978
rect 101318 244294 101374 244350
rect 101442 244294 101498 244350
rect 101318 244170 101374 244226
rect 101442 244170 101498 244226
rect 101318 244046 101374 244102
rect 101442 244046 101498 244102
rect 101318 243922 101374 243978
rect 101442 243922 101498 243978
rect 132038 244294 132094 244350
rect 132162 244294 132218 244350
rect 132038 244170 132094 244226
rect 132162 244170 132218 244226
rect 132038 244046 132094 244102
rect 132162 244046 132218 244102
rect 132038 243922 132094 243978
rect 132162 243922 132218 243978
rect 162758 244294 162814 244350
rect 162882 244294 162938 244350
rect 162758 244170 162814 244226
rect 162882 244170 162938 244226
rect 162758 244046 162814 244102
rect 162882 244046 162938 244102
rect 162758 243922 162814 243978
rect 162882 243922 162938 243978
rect 193478 244294 193534 244350
rect 193602 244294 193658 244350
rect 193478 244170 193534 244226
rect 193602 244170 193658 244226
rect 193478 244046 193534 244102
rect 193602 244046 193658 244102
rect 193478 243922 193534 243978
rect 193602 243922 193658 243978
rect 224198 244294 224254 244350
rect 224322 244294 224378 244350
rect 224198 244170 224254 244226
rect 224322 244170 224378 244226
rect 224198 244046 224254 244102
rect 224322 244046 224378 244102
rect 224198 243922 224254 243978
rect 224322 243922 224378 243978
rect 254918 244294 254974 244350
rect 255042 244294 255098 244350
rect 254918 244170 254974 244226
rect 255042 244170 255098 244226
rect 254918 244046 254974 244102
rect 255042 244046 255098 244102
rect 254918 243922 254974 243978
rect 255042 243922 255098 243978
rect 285638 244294 285694 244350
rect 285762 244294 285818 244350
rect 285638 244170 285694 244226
rect 285762 244170 285818 244226
rect 285638 244046 285694 244102
rect 285762 244046 285818 244102
rect 285638 243922 285694 243978
rect 285762 243922 285818 243978
rect 316358 244294 316414 244350
rect 316482 244294 316538 244350
rect 316358 244170 316414 244226
rect 316482 244170 316538 244226
rect 316358 244046 316414 244102
rect 316482 244046 316538 244102
rect 316358 243922 316414 243978
rect 316482 243922 316538 243978
rect 347078 244294 347134 244350
rect 347202 244294 347258 244350
rect 347078 244170 347134 244226
rect 347202 244170 347258 244226
rect 347078 244046 347134 244102
rect 347202 244046 347258 244102
rect 347078 243922 347134 243978
rect 347202 243922 347258 243978
rect 377798 244294 377854 244350
rect 377922 244294 377978 244350
rect 377798 244170 377854 244226
rect 377922 244170 377978 244226
rect 377798 244046 377854 244102
rect 377922 244046 377978 244102
rect 377798 243922 377854 243978
rect 377922 243922 377978 243978
rect 408518 244294 408574 244350
rect 408642 244294 408698 244350
rect 408518 244170 408574 244226
rect 408642 244170 408698 244226
rect 408518 244046 408574 244102
rect 408642 244046 408698 244102
rect 408518 243922 408574 243978
rect 408642 243922 408698 243978
rect 439238 244294 439294 244350
rect 439362 244294 439418 244350
rect 439238 244170 439294 244226
rect 439362 244170 439418 244226
rect 439238 244046 439294 244102
rect 439362 244046 439418 244102
rect 439238 243922 439294 243978
rect 439362 243922 439418 243978
rect 469958 244294 470014 244350
rect 470082 244294 470138 244350
rect 469958 244170 470014 244226
rect 470082 244170 470138 244226
rect 469958 244046 470014 244102
rect 470082 244046 470138 244102
rect 469958 243922 470014 243978
rect 470082 243922 470138 243978
rect 500678 244294 500734 244350
rect 500802 244294 500858 244350
rect 500678 244170 500734 244226
rect 500802 244170 500858 244226
rect 500678 244046 500734 244102
rect 500802 244046 500858 244102
rect 500678 243922 500734 243978
rect 500802 243922 500858 243978
rect 24518 238294 24574 238350
rect 24642 238294 24698 238350
rect 24518 238170 24574 238226
rect 24642 238170 24698 238226
rect 24518 238046 24574 238102
rect 24642 238046 24698 238102
rect 24518 237922 24574 237978
rect 24642 237922 24698 237978
rect 55238 238294 55294 238350
rect 55362 238294 55418 238350
rect 55238 238170 55294 238226
rect 55362 238170 55418 238226
rect 55238 238046 55294 238102
rect 55362 238046 55418 238102
rect 55238 237922 55294 237978
rect 55362 237922 55418 237978
rect 85958 238294 86014 238350
rect 86082 238294 86138 238350
rect 85958 238170 86014 238226
rect 86082 238170 86138 238226
rect 85958 238046 86014 238102
rect 86082 238046 86138 238102
rect 85958 237922 86014 237978
rect 86082 237922 86138 237978
rect 116678 238294 116734 238350
rect 116802 238294 116858 238350
rect 116678 238170 116734 238226
rect 116802 238170 116858 238226
rect 116678 238046 116734 238102
rect 116802 238046 116858 238102
rect 116678 237922 116734 237978
rect 116802 237922 116858 237978
rect 147398 238294 147454 238350
rect 147522 238294 147578 238350
rect 147398 238170 147454 238226
rect 147522 238170 147578 238226
rect 147398 238046 147454 238102
rect 147522 238046 147578 238102
rect 147398 237922 147454 237978
rect 147522 237922 147578 237978
rect 178118 238294 178174 238350
rect 178242 238294 178298 238350
rect 178118 238170 178174 238226
rect 178242 238170 178298 238226
rect 178118 238046 178174 238102
rect 178242 238046 178298 238102
rect 178118 237922 178174 237978
rect 178242 237922 178298 237978
rect 208838 238294 208894 238350
rect 208962 238294 209018 238350
rect 208838 238170 208894 238226
rect 208962 238170 209018 238226
rect 208838 238046 208894 238102
rect 208962 238046 209018 238102
rect 208838 237922 208894 237978
rect 208962 237922 209018 237978
rect 239558 238294 239614 238350
rect 239682 238294 239738 238350
rect 239558 238170 239614 238226
rect 239682 238170 239738 238226
rect 239558 238046 239614 238102
rect 239682 238046 239738 238102
rect 239558 237922 239614 237978
rect 239682 237922 239738 237978
rect 270278 238294 270334 238350
rect 270402 238294 270458 238350
rect 270278 238170 270334 238226
rect 270402 238170 270458 238226
rect 270278 238046 270334 238102
rect 270402 238046 270458 238102
rect 270278 237922 270334 237978
rect 270402 237922 270458 237978
rect 300998 238294 301054 238350
rect 301122 238294 301178 238350
rect 300998 238170 301054 238226
rect 301122 238170 301178 238226
rect 300998 238046 301054 238102
rect 301122 238046 301178 238102
rect 300998 237922 301054 237978
rect 301122 237922 301178 237978
rect 331718 238294 331774 238350
rect 331842 238294 331898 238350
rect 331718 238170 331774 238226
rect 331842 238170 331898 238226
rect 331718 238046 331774 238102
rect 331842 238046 331898 238102
rect 331718 237922 331774 237978
rect 331842 237922 331898 237978
rect 362438 238294 362494 238350
rect 362562 238294 362618 238350
rect 362438 238170 362494 238226
rect 362562 238170 362618 238226
rect 362438 238046 362494 238102
rect 362562 238046 362618 238102
rect 362438 237922 362494 237978
rect 362562 237922 362618 237978
rect 393158 238294 393214 238350
rect 393282 238294 393338 238350
rect 393158 238170 393214 238226
rect 393282 238170 393338 238226
rect 393158 238046 393214 238102
rect 393282 238046 393338 238102
rect 393158 237922 393214 237978
rect 393282 237922 393338 237978
rect 423878 238294 423934 238350
rect 424002 238294 424058 238350
rect 423878 238170 423934 238226
rect 424002 238170 424058 238226
rect 423878 238046 423934 238102
rect 424002 238046 424058 238102
rect 423878 237922 423934 237978
rect 424002 237922 424058 237978
rect 454598 238294 454654 238350
rect 454722 238294 454778 238350
rect 454598 238170 454654 238226
rect 454722 238170 454778 238226
rect 454598 238046 454654 238102
rect 454722 238046 454778 238102
rect 454598 237922 454654 237978
rect 454722 237922 454778 237978
rect 485318 238294 485374 238350
rect 485442 238294 485498 238350
rect 485318 238170 485374 238226
rect 485442 238170 485498 238226
rect 485318 238046 485374 238102
rect 485442 238046 485498 238102
rect 485318 237922 485374 237978
rect 485442 237922 485498 237978
rect 516038 238294 516094 238350
rect 516162 238294 516218 238350
rect 516038 238170 516094 238226
rect 516162 238170 516218 238226
rect 516038 238046 516094 238102
rect 516162 238046 516218 238102
rect 516038 237922 516094 237978
rect 516162 237922 516218 237978
rect 525250 238294 525306 238350
rect 525374 238294 525430 238350
rect 525498 238294 525554 238350
rect 525622 238294 525678 238350
rect 525250 238170 525306 238226
rect 525374 238170 525430 238226
rect 525498 238170 525554 238226
rect 525622 238170 525678 238226
rect 525250 238046 525306 238102
rect 525374 238046 525430 238102
rect 525498 238046 525554 238102
rect 525622 238046 525678 238102
rect 525250 237922 525306 237978
rect 525374 237922 525430 237978
rect 525498 237922 525554 237978
rect 525622 237922 525678 237978
rect 6970 226294 7026 226350
rect 7094 226294 7150 226350
rect 7218 226294 7274 226350
rect 7342 226294 7398 226350
rect 6970 226170 7026 226226
rect 7094 226170 7150 226226
rect 7218 226170 7274 226226
rect 7342 226170 7398 226226
rect 6970 226046 7026 226102
rect 7094 226046 7150 226102
rect 7218 226046 7274 226102
rect 7342 226046 7398 226102
rect 6970 225922 7026 225978
rect 7094 225922 7150 225978
rect 7218 225922 7274 225978
rect 7342 225922 7398 225978
rect 39878 226294 39934 226350
rect 40002 226294 40058 226350
rect 39878 226170 39934 226226
rect 40002 226170 40058 226226
rect 39878 226046 39934 226102
rect 40002 226046 40058 226102
rect 39878 225922 39934 225978
rect 40002 225922 40058 225978
rect 70598 226294 70654 226350
rect 70722 226294 70778 226350
rect 70598 226170 70654 226226
rect 70722 226170 70778 226226
rect 70598 226046 70654 226102
rect 70722 226046 70778 226102
rect 70598 225922 70654 225978
rect 70722 225922 70778 225978
rect 101318 226294 101374 226350
rect 101442 226294 101498 226350
rect 101318 226170 101374 226226
rect 101442 226170 101498 226226
rect 101318 226046 101374 226102
rect 101442 226046 101498 226102
rect 101318 225922 101374 225978
rect 101442 225922 101498 225978
rect 132038 226294 132094 226350
rect 132162 226294 132218 226350
rect 132038 226170 132094 226226
rect 132162 226170 132218 226226
rect 132038 226046 132094 226102
rect 132162 226046 132218 226102
rect 132038 225922 132094 225978
rect 132162 225922 132218 225978
rect 162758 226294 162814 226350
rect 162882 226294 162938 226350
rect 162758 226170 162814 226226
rect 162882 226170 162938 226226
rect 162758 226046 162814 226102
rect 162882 226046 162938 226102
rect 162758 225922 162814 225978
rect 162882 225922 162938 225978
rect 193478 226294 193534 226350
rect 193602 226294 193658 226350
rect 193478 226170 193534 226226
rect 193602 226170 193658 226226
rect 193478 226046 193534 226102
rect 193602 226046 193658 226102
rect 193478 225922 193534 225978
rect 193602 225922 193658 225978
rect 224198 226294 224254 226350
rect 224322 226294 224378 226350
rect 224198 226170 224254 226226
rect 224322 226170 224378 226226
rect 224198 226046 224254 226102
rect 224322 226046 224378 226102
rect 224198 225922 224254 225978
rect 224322 225922 224378 225978
rect 254918 226294 254974 226350
rect 255042 226294 255098 226350
rect 254918 226170 254974 226226
rect 255042 226170 255098 226226
rect 254918 226046 254974 226102
rect 255042 226046 255098 226102
rect 254918 225922 254974 225978
rect 255042 225922 255098 225978
rect 285638 226294 285694 226350
rect 285762 226294 285818 226350
rect 285638 226170 285694 226226
rect 285762 226170 285818 226226
rect 285638 226046 285694 226102
rect 285762 226046 285818 226102
rect 285638 225922 285694 225978
rect 285762 225922 285818 225978
rect 316358 226294 316414 226350
rect 316482 226294 316538 226350
rect 316358 226170 316414 226226
rect 316482 226170 316538 226226
rect 316358 226046 316414 226102
rect 316482 226046 316538 226102
rect 316358 225922 316414 225978
rect 316482 225922 316538 225978
rect 347078 226294 347134 226350
rect 347202 226294 347258 226350
rect 347078 226170 347134 226226
rect 347202 226170 347258 226226
rect 347078 226046 347134 226102
rect 347202 226046 347258 226102
rect 347078 225922 347134 225978
rect 347202 225922 347258 225978
rect 377798 226294 377854 226350
rect 377922 226294 377978 226350
rect 377798 226170 377854 226226
rect 377922 226170 377978 226226
rect 377798 226046 377854 226102
rect 377922 226046 377978 226102
rect 377798 225922 377854 225978
rect 377922 225922 377978 225978
rect 408518 226294 408574 226350
rect 408642 226294 408698 226350
rect 408518 226170 408574 226226
rect 408642 226170 408698 226226
rect 408518 226046 408574 226102
rect 408642 226046 408698 226102
rect 408518 225922 408574 225978
rect 408642 225922 408698 225978
rect 439238 226294 439294 226350
rect 439362 226294 439418 226350
rect 439238 226170 439294 226226
rect 439362 226170 439418 226226
rect 439238 226046 439294 226102
rect 439362 226046 439418 226102
rect 439238 225922 439294 225978
rect 439362 225922 439418 225978
rect 469958 226294 470014 226350
rect 470082 226294 470138 226350
rect 469958 226170 470014 226226
rect 470082 226170 470138 226226
rect 469958 226046 470014 226102
rect 470082 226046 470138 226102
rect 469958 225922 470014 225978
rect 470082 225922 470138 225978
rect 500678 226294 500734 226350
rect 500802 226294 500858 226350
rect 500678 226170 500734 226226
rect 500802 226170 500858 226226
rect 500678 226046 500734 226102
rect 500802 226046 500858 226102
rect 500678 225922 500734 225978
rect 500802 225922 500858 225978
rect 24518 220294 24574 220350
rect 24642 220294 24698 220350
rect 24518 220170 24574 220226
rect 24642 220170 24698 220226
rect 24518 220046 24574 220102
rect 24642 220046 24698 220102
rect 24518 219922 24574 219978
rect 24642 219922 24698 219978
rect 55238 220294 55294 220350
rect 55362 220294 55418 220350
rect 55238 220170 55294 220226
rect 55362 220170 55418 220226
rect 55238 220046 55294 220102
rect 55362 220046 55418 220102
rect 55238 219922 55294 219978
rect 55362 219922 55418 219978
rect 85958 220294 86014 220350
rect 86082 220294 86138 220350
rect 85958 220170 86014 220226
rect 86082 220170 86138 220226
rect 85958 220046 86014 220102
rect 86082 220046 86138 220102
rect 85958 219922 86014 219978
rect 86082 219922 86138 219978
rect 116678 220294 116734 220350
rect 116802 220294 116858 220350
rect 116678 220170 116734 220226
rect 116802 220170 116858 220226
rect 116678 220046 116734 220102
rect 116802 220046 116858 220102
rect 116678 219922 116734 219978
rect 116802 219922 116858 219978
rect 147398 220294 147454 220350
rect 147522 220294 147578 220350
rect 147398 220170 147454 220226
rect 147522 220170 147578 220226
rect 147398 220046 147454 220102
rect 147522 220046 147578 220102
rect 147398 219922 147454 219978
rect 147522 219922 147578 219978
rect 178118 220294 178174 220350
rect 178242 220294 178298 220350
rect 178118 220170 178174 220226
rect 178242 220170 178298 220226
rect 178118 220046 178174 220102
rect 178242 220046 178298 220102
rect 178118 219922 178174 219978
rect 178242 219922 178298 219978
rect 208838 220294 208894 220350
rect 208962 220294 209018 220350
rect 208838 220170 208894 220226
rect 208962 220170 209018 220226
rect 208838 220046 208894 220102
rect 208962 220046 209018 220102
rect 208838 219922 208894 219978
rect 208962 219922 209018 219978
rect 239558 220294 239614 220350
rect 239682 220294 239738 220350
rect 239558 220170 239614 220226
rect 239682 220170 239738 220226
rect 239558 220046 239614 220102
rect 239682 220046 239738 220102
rect 239558 219922 239614 219978
rect 239682 219922 239738 219978
rect 270278 220294 270334 220350
rect 270402 220294 270458 220350
rect 270278 220170 270334 220226
rect 270402 220170 270458 220226
rect 270278 220046 270334 220102
rect 270402 220046 270458 220102
rect 270278 219922 270334 219978
rect 270402 219922 270458 219978
rect 300998 220294 301054 220350
rect 301122 220294 301178 220350
rect 300998 220170 301054 220226
rect 301122 220170 301178 220226
rect 300998 220046 301054 220102
rect 301122 220046 301178 220102
rect 300998 219922 301054 219978
rect 301122 219922 301178 219978
rect 331718 220294 331774 220350
rect 331842 220294 331898 220350
rect 331718 220170 331774 220226
rect 331842 220170 331898 220226
rect 331718 220046 331774 220102
rect 331842 220046 331898 220102
rect 331718 219922 331774 219978
rect 331842 219922 331898 219978
rect 362438 220294 362494 220350
rect 362562 220294 362618 220350
rect 362438 220170 362494 220226
rect 362562 220170 362618 220226
rect 362438 220046 362494 220102
rect 362562 220046 362618 220102
rect 362438 219922 362494 219978
rect 362562 219922 362618 219978
rect 393158 220294 393214 220350
rect 393282 220294 393338 220350
rect 393158 220170 393214 220226
rect 393282 220170 393338 220226
rect 393158 220046 393214 220102
rect 393282 220046 393338 220102
rect 393158 219922 393214 219978
rect 393282 219922 393338 219978
rect 423878 220294 423934 220350
rect 424002 220294 424058 220350
rect 423878 220170 423934 220226
rect 424002 220170 424058 220226
rect 423878 220046 423934 220102
rect 424002 220046 424058 220102
rect 423878 219922 423934 219978
rect 424002 219922 424058 219978
rect 454598 220294 454654 220350
rect 454722 220294 454778 220350
rect 454598 220170 454654 220226
rect 454722 220170 454778 220226
rect 454598 220046 454654 220102
rect 454722 220046 454778 220102
rect 454598 219922 454654 219978
rect 454722 219922 454778 219978
rect 485318 220294 485374 220350
rect 485442 220294 485498 220350
rect 485318 220170 485374 220226
rect 485442 220170 485498 220226
rect 485318 220046 485374 220102
rect 485442 220046 485498 220102
rect 485318 219922 485374 219978
rect 485442 219922 485498 219978
rect 516038 220294 516094 220350
rect 516162 220294 516218 220350
rect 516038 220170 516094 220226
rect 516162 220170 516218 220226
rect 516038 220046 516094 220102
rect 516162 220046 516218 220102
rect 516038 219922 516094 219978
rect 516162 219922 516218 219978
rect 525250 220294 525306 220350
rect 525374 220294 525430 220350
rect 525498 220294 525554 220350
rect 525622 220294 525678 220350
rect 525250 220170 525306 220226
rect 525374 220170 525430 220226
rect 525498 220170 525554 220226
rect 525622 220170 525678 220226
rect 525250 220046 525306 220102
rect 525374 220046 525430 220102
rect 525498 220046 525554 220102
rect 525622 220046 525678 220102
rect 525250 219922 525306 219978
rect 525374 219922 525430 219978
rect 525498 219922 525554 219978
rect 525622 219922 525678 219978
rect 6970 208294 7026 208350
rect 7094 208294 7150 208350
rect 7218 208294 7274 208350
rect 7342 208294 7398 208350
rect 6970 208170 7026 208226
rect 7094 208170 7150 208226
rect 7218 208170 7274 208226
rect 7342 208170 7398 208226
rect 6970 208046 7026 208102
rect 7094 208046 7150 208102
rect 7218 208046 7274 208102
rect 7342 208046 7398 208102
rect 6970 207922 7026 207978
rect 7094 207922 7150 207978
rect 7218 207922 7274 207978
rect 7342 207922 7398 207978
rect 39878 208294 39934 208350
rect 40002 208294 40058 208350
rect 39878 208170 39934 208226
rect 40002 208170 40058 208226
rect 39878 208046 39934 208102
rect 40002 208046 40058 208102
rect 39878 207922 39934 207978
rect 40002 207922 40058 207978
rect 70598 208294 70654 208350
rect 70722 208294 70778 208350
rect 70598 208170 70654 208226
rect 70722 208170 70778 208226
rect 70598 208046 70654 208102
rect 70722 208046 70778 208102
rect 70598 207922 70654 207978
rect 70722 207922 70778 207978
rect 101318 208294 101374 208350
rect 101442 208294 101498 208350
rect 101318 208170 101374 208226
rect 101442 208170 101498 208226
rect 101318 208046 101374 208102
rect 101442 208046 101498 208102
rect 101318 207922 101374 207978
rect 101442 207922 101498 207978
rect 132038 208294 132094 208350
rect 132162 208294 132218 208350
rect 132038 208170 132094 208226
rect 132162 208170 132218 208226
rect 132038 208046 132094 208102
rect 132162 208046 132218 208102
rect 132038 207922 132094 207978
rect 132162 207922 132218 207978
rect 162758 208294 162814 208350
rect 162882 208294 162938 208350
rect 162758 208170 162814 208226
rect 162882 208170 162938 208226
rect 162758 208046 162814 208102
rect 162882 208046 162938 208102
rect 162758 207922 162814 207978
rect 162882 207922 162938 207978
rect 193478 208294 193534 208350
rect 193602 208294 193658 208350
rect 193478 208170 193534 208226
rect 193602 208170 193658 208226
rect 193478 208046 193534 208102
rect 193602 208046 193658 208102
rect 193478 207922 193534 207978
rect 193602 207922 193658 207978
rect 224198 208294 224254 208350
rect 224322 208294 224378 208350
rect 224198 208170 224254 208226
rect 224322 208170 224378 208226
rect 224198 208046 224254 208102
rect 224322 208046 224378 208102
rect 224198 207922 224254 207978
rect 224322 207922 224378 207978
rect 254918 208294 254974 208350
rect 255042 208294 255098 208350
rect 254918 208170 254974 208226
rect 255042 208170 255098 208226
rect 254918 208046 254974 208102
rect 255042 208046 255098 208102
rect 254918 207922 254974 207978
rect 255042 207922 255098 207978
rect 285638 208294 285694 208350
rect 285762 208294 285818 208350
rect 285638 208170 285694 208226
rect 285762 208170 285818 208226
rect 285638 208046 285694 208102
rect 285762 208046 285818 208102
rect 285638 207922 285694 207978
rect 285762 207922 285818 207978
rect 316358 208294 316414 208350
rect 316482 208294 316538 208350
rect 316358 208170 316414 208226
rect 316482 208170 316538 208226
rect 316358 208046 316414 208102
rect 316482 208046 316538 208102
rect 316358 207922 316414 207978
rect 316482 207922 316538 207978
rect 347078 208294 347134 208350
rect 347202 208294 347258 208350
rect 347078 208170 347134 208226
rect 347202 208170 347258 208226
rect 347078 208046 347134 208102
rect 347202 208046 347258 208102
rect 347078 207922 347134 207978
rect 347202 207922 347258 207978
rect 377798 208294 377854 208350
rect 377922 208294 377978 208350
rect 377798 208170 377854 208226
rect 377922 208170 377978 208226
rect 377798 208046 377854 208102
rect 377922 208046 377978 208102
rect 377798 207922 377854 207978
rect 377922 207922 377978 207978
rect 408518 208294 408574 208350
rect 408642 208294 408698 208350
rect 408518 208170 408574 208226
rect 408642 208170 408698 208226
rect 408518 208046 408574 208102
rect 408642 208046 408698 208102
rect 408518 207922 408574 207978
rect 408642 207922 408698 207978
rect 439238 208294 439294 208350
rect 439362 208294 439418 208350
rect 439238 208170 439294 208226
rect 439362 208170 439418 208226
rect 439238 208046 439294 208102
rect 439362 208046 439418 208102
rect 439238 207922 439294 207978
rect 439362 207922 439418 207978
rect 469958 208294 470014 208350
rect 470082 208294 470138 208350
rect 469958 208170 470014 208226
rect 470082 208170 470138 208226
rect 469958 208046 470014 208102
rect 470082 208046 470138 208102
rect 469958 207922 470014 207978
rect 470082 207922 470138 207978
rect 500678 208294 500734 208350
rect 500802 208294 500858 208350
rect 500678 208170 500734 208226
rect 500802 208170 500858 208226
rect 500678 208046 500734 208102
rect 500802 208046 500858 208102
rect 500678 207922 500734 207978
rect 500802 207922 500858 207978
rect 24518 202294 24574 202350
rect 24642 202294 24698 202350
rect 24518 202170 24574 202226
rect 24642 202170 24698 202226
rect 24518 202046 24574 202102
rect 24642 202046 24698 202102
rect 24518 201922 24574 201978
rect 24642 201922 24698 201978
rect 55238 202294 55294 202350
rect 55362 202294 55418 202350
rect 55238 202170 55294 202226
rect 55362 202170 55418 202226
rect 55238 202046 55294 202102
rect 55362 202046 55418 202102
rect 55238 201922 55294 201978
rect 55362 201922 55418 201978
rect 85958 202294 86014 202350
rect 86082 202294 86138 202350
rect 85958 202170 86014 202226
rect 86082 202170 86138 202226
rect 85958 202046 86014 202102
rect 86082 202046 86138 202102
rect 85958 201922 86014 201978
rect 86082 201922 86138 201978
rect 116678 202294 116734 202350
rect 116802 202294 116858 202350
rect 116678 202170 116734 202226
rect 116802 202170 116858 202226
rect 116678 202046 116734 202102
rect 116802 202046 116858 202102
rect 116678 201922 116734 201978
rect 116802 201922 116858 201978
rect 147398 202294 147454 202350
rect 147522 202294 147578 202350
rect 147398 202170 147454 202226
rect 147522 202170 147578 202226
rect 147398 202046 147454 202102
rect 147522 202046 147578 202102
rect 147398 201922 147454 201978
rect 147522 201922 147578 201978
rect 178118 202294 178174 202350
rect 178242 202294 178298 202350
rect 178118 202170 178174 202226
rect 178242 202170 178298 202226
rect 178118 202046 178174 202102
rect 178242 202046 178298 202102
rect 178118 201922 178174 201978
rect 178242 201922 178298 201978
rect 208838 202294 208894 202350
rect 208962 202294 209018 202350
rect 208838 202170 208894 202226
rect 208962 202170 209018 202226
rect 208838 202046 208894 202102
rect 208962 202046 209018 202102
rect 208838 201922 208894 201978
rect 208962 201922 209018 201978
rect 239558 202294 239614 202350
rect 239682 202294 239738 202350
rect 239558 202170 239614 202226
rect 239682 202170 239738 202226
rect 239558 202046 239614 202102
rect 239682 202046 239738 202102
rect 239558 201922 239614 201978
rect 239682 201922 239738 201978
rect 270278 202294 270334 202350
rect 270402 202294 270458 202350
rect 270278 202170 270334 202226
rect 270402 202170 270458 202226
rect 270278 202046 270334 202102
rect 270402 202046 270458 202102
rect 270278 201922 270334 201978
rect 270402 201922 270458 201978
rect 300998 202294 301054 202350
rect 301122 202294 301178 202350
rect 300998 202170 301054 202226
rect 301122 202170 301178 202226
rect 300998 202046 301054 202102
rect 301122 202046 301178 202102
rect 300998 201922 301054 201978
rect 301122 201922 301178 201978
rect 331718 202294 331774 202350
rect 331842 202294 331898 202350
rect 331718 202170 331774 202226
rect 331842 202170 331898 202226
rect 331718 202046 331774 202102
rect 331842 202046 331898 202102
rect 331718 201922 331774 201978
rect 331842 201922 331898 201978
rect 362438 202294 362494 202350
rect 362562 202294 362618 202350
rect 362438 202170 362494 202226
rect 362562 202170 362618 202226
rect 362438 202046 362494 202102
rect 362562 202046 362618 202102
rect 362438 201922 362494 201978
rect 362562 201922 362618 201978
rect 393158 202294 393214 202350
rect 393282 202294 393338 202350
rect 393158 202170 393214 202226
rect 393282 202170 393338 202226
rect 393158 202046 393214 202102
rect 393282 202046 393338 202102
rect 393158 201922 393214 201978
rect 393282 201922 393338 201978
rect 423878 202294 423934 202350
rect 424002 202294 424058 202350
rect 423878 202170 423934 202226
rect 424002 202170 424058 202226
rect 423878 202046 423934 202102
rect 424002 202046 424058 202102
rect 423878 201922 423934 201978
rect 424002 201922 424058 201978
rect 454598 202294 454654 202350
rect 454722 202294 454778 202350
rect 454598 202170 454654 202226
rect 454722 202170 454778 202226
rect 454598 202046 454654 202102
rect 454722 202046 454778 202102
rect 454598 201922 454654 201978
rect 454722 201922 454778 201978
rect 485318 202294 485374 202350
rect 485442 202294 485498 202350
rect 485318 202170 485374 202226
rect 485442 202170 485498 202226
rect 485318 202046 485374 202102
rect 485442 202046 485498 202102
rect 485318 201922 485374 201978
rect 485442 201922 485498 201978
rect 516038 202294 516094 202350
rect 516162 202294 516218 202350
rect 516038 202170 516094 202226
rect 516162 202170 516218 202226
rect 516038 202046 516094 202102
rect 516162 202046 516218 202102
rect 516038 201922 516094 201978
rect 516162 201922 516218 201978
rect 525250 202294 525306 202350
rect 525374 202294 525430 202350
rect 525498 202294 525554 202350
rect 525622 202294 525678 202350
rect 525250 202170 525306 202226
rect 525374 202170 525430 202226
rect 525498 202170 525554 202226
rect 525622 202170 525678 202226
rect 525250 202046 525306 202102
rect 525374 202046 525430 202102
rect 525498 202046 525554 202102
rect 525622 202046 525678 202102
rect 525250 201922 525306 201978
rect 525374 201922 525430 201978
rect 525498 201922 525554 201978
rect 525622 201922 525678 201978
rect 6970 190294 7026 190350
rect 7094 190294 7150 190350
rect 7218 190294 7274 190350
rect 7342 190294 7398 190350
rect 6970 190170 7026 190226
rect 7094 190170 7150 190226
rect 7218 190170 7274 190226
rect 7342 190170 7398 190226
rect 6970 190046 7026 190102
rect 7094 190046 7150 190102
rect 7218 190046 7274 190102
rect 7342 190046 7398 190102
rect 6970 189922 7026 189978
rect 7094 189922 7150 189978
rect 7218 189922 7274 189978
rect 7342 189922 7398 189978
rect 39878 190294 39934 190350
rect 40002 190294 40058 190350
rect 39878 190170 39934 190226
rect 40002 190170 40058 190226
rect 39878 190046 39934 190102
rect 40002 190046 40058 190102
rect 39878 189922 39934 189978
rect 40002 189922 40058 189978
rect 70598 190294 70654 190350
rect 70722 190294 70778 190350
rect 70598 190170 70654 190226
rect 70722 190170 70778 190226
rect 70598 190046 70654 190102
rect 70722 190046 70778 190102
rect 70598 189922 70654 189978
rect 70722 189922 70778 189978
rect 101318 190294 101374 190350
rect 101442 190294 101498 190350
rect 101318 190170 101374 190226
rect 101442 190170 101498 190226
rect 101318 190046 101374 190102
rect 101442 190046 101498 190102
rect 101318 189922 101374 189978
rect 101442 189922 101498 189978
rect 132038 190294 132094 190350
rect 132162 190294 132218 190350
rect 132038 190170 132094 190226
rect 132162 190170 132218 190226
rect 132038 190046 132094 190102
rect 132162 190046 132218 190102
rect 132038 189922 132094 189978
rect 132162 189922 132218 189978
rect 162758 190294 162814 190350
rect 162882 190294 162938 190350
rect 162758 190170 162814 190226
rect 162882 190170 162938 190226
rect 162758 190046 162814 190102
rect 162882 190046 162938 190102
rect 162758 189922 162814 189978
rect 162882 189922 162938 189978
rect 193478 190294 193534 190350
rect 193602 190294 193658 190350
rect 193478 190170 193534 190226
rect 193602 190170 193658 190226
rect 193478 190046 193534 190102
rect 193602 190046 193658 190102
rect 193478 189922 193534 189978
rect 193602 189922 193658 189978
rect 224198 190294 224254 190350
rect 224322 190294 224378 190350
rect 224198 190170 224254 190226
rect 224322 190170 224378 190226
rect 224198 190046 224254 190102
rect 224322 190046 224378 190102
rect 224198 189922 224254 189978
rect 224322 189922 224378 189978
rect 254918 190294 254974 190350
rect 255042 190294 255098 190350
rect 254918 190170 254974 190226
rect 255042 190170 255098 190226
rect 254918 190046 254974 190102
rect 255042 190046 255098 190102
rect 254918 189922 254974 189978
rect 255042 189922 255098 189978
rect 285638 190294 285694 190350
rect 285762 190294 285818 190350
rect 285638 190170 285694 190226
rect 285762 190170 285818 190226
rect 285638 190046 285694 190102
rect 285762 190046 285818 190102
rect 285638 189922 285694 189978
rect 285762 189922 285818 189978
rect 316358 190294 316414 190350
rect 316482 190294 316538 190350
rect 316358 190170 316414 190226
rect 316482 190170 316538 190226
rect 316358 190046 316414 190102
rect 316482 190046 316538 190102
rect 316358 189922 316414 189978
rect 316482 189922 316538 189978
rect 347078 190294 347134 190350
rect 347202 190294 347258 190350
rect 347078 190170 347134 190226
rect 347202 190170 347258 190226
rect 347078 190046 347134 190102
rect 347202 190046 347258 190102
rect 347078 189922 347134 189978
rect 347202 189922 347258 189978
rect 377798 190294 377854 190350
rect 377922 190294 377978 190350
rect 377798 190170 377854 190226
rect 377922 190170 377978 190226
rect 377798 190046 377854 190102
rect 377922 190046 377978 190102
rect 377798 189922 377854 189978
rect 377922 189922 377978 189978
rect 408518 190294 408574 190350
rect 408642 190294 408698 190350
rect 408518 190170 408574 190226
rect 408642 190170 408698 190226
rect 408518 190046 408574 190102
rect 408642 190046 408698 190102
rect 408518 189922 408574 189978
rect 408642 189922 408698 189978
rect 439238 190294 439294 190350
rect 439362 190294 439418 190350
rect 439238 190170 439294 190226
rect 439362 190170 439418 190226
rect 439238 190046 439294 190102
rect 439362 190046 439418 190102
rect 439238 189922 439294 189978
rect 439362 189922 439418 189978
rect 469958 190294 470014 190350
rect 470082 190294 470138 190350
rect 469958 190170 470014 190226
rect 470082 190170 470138 190226
rect 469958 190046 470014 190102
rect 470082 190046 470138 190102
rect 469958 189922 470014 189978
rect 470082 189922 470138 189978
rect 500678 190294 500734 190350
rect 500802 190294 500858 190350
rect 500678 190170 500734 190226
rect 500802 190170 500858 190226
rect 500678 190046 500734 190102
rect 500802 190046 500858 190102
rect 500678 189922 500734 189978
rect 500802 189922 500858 189978
rect 24518 184294 24574 184350
rect 24642 184294 24698 184350
rect 24518 184170 24574 184226
rect 24642 184170 24698 184226
rect 24518 184046 24574 184102
rect 24642 184046 24698 184102
rect 24518 183922 24574 183978
rect 24642 183922 24698 183978
rect 55238 184294 55294 184350
rect 55362 184294 55418 184350
rect 55238 184170 55294 184226
rect 55362 184170 55418 184226
rect 55238 184046 55294 184102
rect 55362 184046 55418 184102
rect 55238 183922 55294 183978
rect 55362 183922 55418 183978
rect 85958 184294 86014 184350
rect 86082 184294 86138 184350
rect 85958 184170 86014 184226
rect 86082 184170 86138 184226
rect 85958 184046 86014 184102
rect 86082 184046 86138 184102
rect 85958 183922 86014 183978
rect 86082 183922 86138 183978
rect 116678 184294 116734 184350
rect 116802 184294 116858 184350
rect 116678 184170 116734 184226
rect 116802 184170 116858 184226
rect 116678 184046 116734 184102
rect 116802 184046 116858 184102
rect 116678 183922 116734 183978
rect 116802 183922 116858 183978
rect 147398 184294 147454 184350
rect 147522 184294 147578 184350
rect 147398 184170 147454 184226
rect 147522 184170 147578 184226
rect 147398 184046 147454 184102
rect 147522 184046 147578 184102
rect 147398 183922 147454 183978
rect 147522 183922 147578 183978
rect 178118 184294 178174 184350
rect 178242 184294 178298 184350
rect 178118 184170 178174 184226
rect 178242 184170 178298 184226
rect 178118 184046 178174 184102
rect 178242 184046 178298 184102
rect 178118 183922 178174 183978
rect 178242 183922 178298 183978
rect 208838 184294 208894 184350
rect 208962 184294 209018 184350
rect 208838 184170 208894 184226
rect 208962 184170 209018 184226
rect 208838 184046 208894 184102
rect 208962 184046 209018 184102
rect 208838 183922 208894 183978
rect 208962 183922 209018 183978
rect 239558 184294 239614 184350
rect 239682 184294 239738 184350
rect 239558 184170 239614 184226
rect 239682 184170 239738 184226
rect 239558 184046 239614 184102
rect 239682 184046 239738 184102
rect 239558 183922 239614 183978
rect 239682 183922 239738 183978
rect 270278 184294 270334 184350
rect 270402 184294 270458 184350
rect 270278 184170 270334 184226
rect 270402 184170 270458 184226
rect 270278 184046 270334 184102
rect 270402 184046 270458 184102
rect 270278 183922 270334 183978
rect 270402 183922 270458 183978
rect 300998 184294 301054 184350
rect 301122 184294 301178 184350
rect 300998 184170 301054 184226
rect 301122 184170 301178 184226
rect 300998 184046 301054 184102
rect 301122 184046 301178 184102
rect 300998 183922 301054 183978
rect 301122 183922 301178 183978
rect 331718 184294 331774 184350
rect 331842 184294 331898 184350
rect 331718 184170 331774 184226
rect 331842 184170 331898 184226
rect 331718 184046 331774 184102
rect 331842 184046 331898 184102
rect 331718 183922 331774 183978
rect 331842 183922 331898 183978
rect 362438 184294 362494 184350
rect 362562 184294 362618 184350
rect 362438 184170 362494 184226
rect 362562 184170 362618 184226
rect 362438 184046 362494 184102
rect 362562 184046 362618 184102
rect 362438 183922 362494 183978
rect 362562 183922 362618 183978
rect 393158 184294 393214 184350
rect 393282 184294 393338 184350
rect 393158 184170 393214 184226
rect 393282 184170 393338 184226
rect 393158 184046 393214 184102
rect 393282 184046 393338 184102
rect 393158 183922 393214 183978
rect 393282 183922 393338 183978
rect 423878 184294 423934 184350
rect 424002 184294 424058 184350
rect 423878 184170 423934 184226
rect 424002 184170 424058 184226
rect 423878 184046 423934 184102
rect 424002 184046 424058 184102
rect 423878 183922 423934 183978
rect 424002 183922 424058 183978
rect 454598 184294 454654 184350
rect 454722 184294 454778 184350
rect 454598 184170 454654 184226
rect 454722 184170 454778 184226
rect 454598 184046 454654 184102
rect 454722 184046 454778 184102
rect 454598 183922 454654 183978
rect 454722 183922 454778 183978
rect 485318 184294 485374 184350
rect 485442 184294 485498 184350
rect 485318 184170 485374 184226
rect 485442 184170 485498 184226
rect 485318 184046 485374 184102
rect 485442 184046 485498 184102
rect 485318 183922 485374 183978
rect 485442 183922 485498 183978
rect 516038 184294 516094 184350
rect 516162 184294 516218 184350
rect 516038 184170 516094 184226
rect 516162 184170 516218 184226
rect 516038 184046 516094 184102
rect 516162 184046 516218 184102
rect 516038 183922 516094 183978
rect 516162 183922 516218 183978
rect 525250 184294 525306 184350
rect 525374 184294 525430 184350
rect 525498 184294 525554 184350
rect 525622 184294 525678 184350
rect 525250 184170 525306 184226
rect 525374 184170 525430 184226
rect 525498 184170 525554 184226
rect 525622 184170 525678 184226
rect 525250 184046 525306 184102
rect 525374 184046 525430 184102
rect 525498 184046 525554 184102
rect 525622 184046 525678 184102
rect 525250 183922 525306 183978
rect 525374 183922 525430 183978
rect 525498 183922 525554 183978
rect 525622 183922 525678 183978
rect 6970 172294 7026 172350
rect 7094 172294 7150 172350
rect 7218 172294 7274 172350
rect 7342 172294 7398 172350
rect 6970 172170 7026 172226
rect 7094 172170 7150 172226
rect 7218 172170 7274 172226
rect 7342 172170 7398 172226
rect 6970 172046 7026 172102
rect 7094 172046 7150 172102
rect 7218 172046 7274 172102
rect 7342 172046 7398 172102
rect 6970 171922 7026 171978
rect 7094 171922 7150 171978
rect 7218 171922 7274 171978
rect 7342 171922 7398 171978
rect 39878 172294 39934 172350
rect 40002 172294 40058 172350
rect 39878 172170 39934 172226
rect 40002 172170 40058 172226
rect 39878 172046 39934 172102
rect 40002 172046 40058 172102
rect 39878 171922 39934 171978
rect 40002 171922 40058 171978
rect 70598 172294 70654 172350
rect 70722 172294 70778 172350
rect 70598 172170 70654 172226
rect 70722 172170 70778 172226
rect 70598 172046 70654 172102
rect 70722 172046 70778 172102
rect 70598 171922 70654 171978
rect 70722 171922 70778 171978
rect 101318 172294 101374 172350
rect 101442 172294 101498 172350
rect 101318 172170 101374 172226
rect 101442 172170 101498 172226
rect 101318 172046 101374 172102
rect 101442 172046 101498 172102
rect 101318 171922 101374 171978
rect 101442 171922 101498 171978
rect 132038 172294 132094 172350
rect 132162 172294 132218 172350
rect 132038 172170 132094 172226
rect 132162 172170 132218 172226
rect 132038 172046 132094 172102
rect 132162 172046 132218 172102
rect 132038 171922 132094 171978
rect 132162 171922 132218 171978
rect 162758 172294 162814 172350
rect 162882 172294 162938 172350
rect 162758 172170 162814 172226
rect 162882 172170 162938 172226
rect 162758 172046 162814 172102
rect 162882 172046 162938 172102
rect 162758 171922 162814 171978
rect 162882 171922 162938 171978
rect 193478 172294 193534 172350
rect 193602 172294 193658 172350
rect 193478 172170 193534 172226
rect 193602 172170 193658 172226
rect 193478 172046 193534 172102
rect 193602 172046 193658 172102
rect 193478 171922 193534 171978
rect 193602 171922 193658 171978
rect 224198 172294 224254 172350
rect 224322 172294 224378 172350
rect 224198 172170 224254 172226
rect 224322 172170 224378 172226
rect 224198 172046 224254 172102
rect 224322 172046 224378 172102
rect 224198 171922 224254 171978
rect 224322 171922 224378 171978
rect 254918 172294 254974 172350
rect 255042 172294 255098 172350
rect 254918 172170 254974 172226
rect 255042 172170 255098 172226
rect 254918 172046 254974 172102
rect 255042 172046 255098 172102
rect 254918 171922 254974 171978
rect 255042 171922 255098 171978
rect 285638 172294 285694 172350
rect 285762 172294 285818 172350
rect 285638 172170 285694 172226
rect 285762 172170 285818 172226
rect 285638 172046 285694 172102
rect 285762 172046 285818 172102
rect 285638 171922 285694 171978
rect 285762 171922 285818 171978
rect 316358 172294 316414 172350
rect 316482 172294 316538 172350
rect 316358 172170 316414 172226
rect 316482 172170 316538 172226
rect 316358 172046 316414 172102
rect 316482 172046 316538 172102
rect 316358 171922 316414 171978
rect 316482 171922 316538 171978
rect 347078 172294 347134 172350
rect 347202 172294 347258 172350
rect 347078 172170 347134 172226
rect 347202 172170 347258 172226
rect 347078 172046 347134 172102
rect 347202 172046 347258 172102
rect 347078 171922 347134 171978
rect 347202 171922 347258 171978
rect 377798 172294 377854 172350
rect 377922 172294 377978 172350
rect 377798 172170 377854 172226
rect 377922 172170 377978 172226
rect 377798 172046 377854 172102
rect 377922 172046 377978 172102
rect 377798 171922 377854 171978
rect 377922 171922 377978 171978
rect 408518 172294 408574 172350
rect 408642 172294 408698 172350
rect 408518 172170 408574 172226
rect 408642 172170 408698 172226
rect 408518 172046 408574 172102
rect 408642 172046 408698 172102
rect 408518 171922 408574 171978
rect 408642 171922 408698 171978
rect 439238 172294 439294 172350
rect 439362 172294 439418 172350
rect 439238 172170 439294 172226
rect 439362 172170 439418 172226
rect 439238 172046 439294 172102
rect 439362 172046 439418 172102
rect 439238 171922 439294 171978
rect 439362 171922 439418 171978
rect 469958 172294 470014 172350
rect 470082 172294 470138 172350
rect 469958 172170 470014 172226
rect 470082 172170 470138 172226
rect 469958 172046 470014 172102
rect 470082 172046 470138 172102
rect 469958 171922 470014 171978
rect 470082 171922 470138 171978
rect 500678 172294 500734 172350
rect 500802 172294 500858 172350
rect 500678 172170 500734 172226
rect 500802 172170 500858 172226
rect 500678 172046 500734 172102
rect 500802 172046 500858 172102
rect 500678 171922 500734 171978
rect 500802 171922 500858 171978
rect 24518 166294 24574 166350
rect 24642 166294 24698 166350
rect 24518 166170 24574 166226
rect 24642 166170 24698 166226
rect 24518 166046 24574 166102
rect 24642 166046 24698 166102
rect 24518 165922 24574 165978
rect 24642 165922 24698 165978
rect 55238 166294 55294 166350
rect 55362 166294 55418 166350
rect 55238 166170 55294 166226
rect 55362 166170 55418 166226
rect 55238 166046 55294 166102
rect 55362 166046 55418 166102
rect 55238 165922 55294 165978
rect 55362 165922 55418 165978
rect 85958 166294 86014 166350
rect 86082 166294 86138 166350
rect 85958 166170 86014 166226
rect 86082 166170 86138 166226
rect 85958 166046 86014 166102
rect 86082 166046 86138 166102
rect 85958 165922 86014 165978
rect 86082 165922 86138 165978
rect 116678 166294 116734 166350
rect 116802 166294 116858 166350
rect 116678 166170 116734 166226
rect 116802 166170 116858 166226
rect 116678 166046 116734 166102
rect 116802 166046 116858 166102
rect 116678 165922 116734 165978
rect 116802 165922 116858 165978
rect 147398 166294 147454 166350
rect 147522 166294 147578 166350
rect 147398 166170 147454 166226
rect 147522 166170 147578 166226
rect 147398 166046 147454 166102
rect 147522 166046 147578 166102
rect 147398 165922 147454 165978
rect 147522 165922 147578 165978
rect 178118 166294 178174 166350
rect 178242 166294 178298 166350
rect 178118 166170 178174 166226
rect 178242 166170 178298 166226
rect 178118 166046 178174 166102
rect 178242 166046 178298 166102
rect 178118 165922 178174 165978
rect 178242 165922 178298 165978
rect 208838 166294 208894 166350
rect 208962 166294 209018 166350
rect 208838 166170 208894 166226
rect 208962 166170 209018 166226
rect 208838 166046 208894 166102
rect 208962 166046 209018 166102
rect 208838 165922 208894 165978
rect 208962 165922 209018 165978
rect 239558 166294 239614 166350
rect 239682 166294 239738 166350
rect 239558 166170 239614 166226
rect 239682 166170 239738 166226
rect 239558 166046 239614 166102
rect 239682 166046 239738 166102
rect 239558 165922 239614 165978
rect 239682 165922 239738 165978
rect 270278 166294 270334 166350
rect 270402 166294 270458 166350
rect 270278 166170 270334 166226
rect 270402 166170 270458 166226
rect 270278 166046 270334 166102
rect 270402 166046 270458 166102
rect 270278 165922 270334 165978
rect 270402 165922 270458 165978
rect 300998 166294 301054 166350
rect 301122 166294 301178 166350
rect 300998 166170 301054 166226
rect 301122 166170 301178 166226
rect 300998 166046 301054 166102
rect 301122 166046 301178 166102
rect 300998 165922 301054 165978
rect 301122 165922 301178 165978
rect 331718 166294 331774 166350
rect 331842 166294 331898 166350
rect 331718 166170 331774 166226
rect 331842 166170 331898 166226
rect 331718 166046 331774 166102
rect 331842 166046 331898 166102
rect 331718 165922 331774 165978
rect 331842 165922 331898 165978
rect 362438 166294 362494 166350
rect 362562 166294 362618 166350
rect 362438 166170 362494 166226
rect 362562 166170 362618 166226
rect 362438 166046 362494 166102
rect 362562 166046 362618 166102
rect 362438 165922 362494 165978
rect 362562 165922 362618 165978
rect 393158 166294 393214 166350
rect 393282 166294 393338 166350
rect 393158 166170 393214 166226
rect 393282 166170 393338 166226
rect 393158 166046 393214 166102
rect 393282 166046 393338 166102
rect 393158 165922 393214 165978
rect 393282 165922 393338 165978
rect 423878 166294 423934 166350
rect 424002 166294 424058 166350
rect 423878 166170 423934 166226
rect 424002 166170 424058 166226
rect 423878 166046 423934 166102
rect 424002 166046 424058 166102
rect 423878 165922 423934 165978
rect 424002 165922 424058 165978
rect 454598 166294 454654 166350
rect 454722 166294 454778 166350
rect 454598 166170 454654 166226
rect 454722 166170 454778 166226
rect 454598 166046 454654 166102
rect 454722 166046 454778 166102
rect 454598 165922 454654 165978
rect 454722 165922 454778 165978
rect 485318 166294 485374 166350
rect 485442 166294 485498 166350
rect 485318 166170 485374 166226
rect 485442 166170 485498 166226
rect 485318 166046 485374 166102
rect 485442 166046 485498 166102
rect 485318 165922 485374 165978
rect 485442 165922 485498 165978
rect 516038 166294 516094 166350
rect 516162 166294 516218 166350
rect 516038 166170 516094 166226
rect 516162 166170 516218 166226
rect 516038 166046 516094 166102
rect 516162 166046 516218 166102
rect 516038 165922 516094 165978
rect 516162 165922 516218 165978
rect 525250 166294 525306 166350
rect 525374 166294 525430 166350
rect 525498 166294 525554 166350
rect 525622 166294 525678 166350
rect 525250 166170 525306 166226
rect 525374 166170 525430 166226
rect 525498 166170 525554 166226
rect 525622 166170 525678 166226
rect 525250 166046 525306 166102
rect 525374 166046 525430 166102
rect 525498 166046 525554 166102
rect 525622 166046 525678 166102
rect 525250 165922 525306 165978
rect 525374 165922 525430 165978
rect 525498 165922 525554 165978
rect 525622 165922 525678 165978
rect 6970 154294 7026 154350
rect 7094 154294 7150 154350
rect 7218 154294 7274 154350
rect 7342 154294 7398 154350
rect 6970 154170 7026 154226
rect 7094 154170 7150 154226
rect 7218 154170 7274 154226
rect 7342 154170 7398 154226
rect 6970 154046 7026 154102
rect 7094 154046 7150 154102
rect 7218 154046 7274 154102
rect 7342 154046 7398 154102
rect 6970 153922 7026 153978
rect 7094 153922 7150 153978
rect 7218 153922 7274 153978
rect 7342 153922 7398 153978
rect 39878 154294 39934 154350
rect 40002 154294 40058 154350
rect 39878 154170 39934 154226
rect 40002 154170 40058 154226
rect 39878 154046 39934 154102
rect 40002 154046 40058 154102
rect 39878 153922 39934 153978
rect 40002 153922 40058 153978
rect 70598 154294 70654 154350
rect 70722 154294 70778 154350
rect 70598 154170 70654 154226
rect 70722 154170 70778 154226
rect 70598 154046 70654 154102
rect 70722 154046 70778 154102
rect 70598 153922 70654 153978
rect 70722 153922 70778 153978
rect 101318 154294 101374 154350
rect 101442 154294 101498 154350
rect 101318 154170 101374 154226
rect 101442 154170 101498 154226
rect 101318 154046 101374 154102
rect 101442 154046 101498 154102
rect 101318 153922 101374 153978
rect 101442 153922 101498 153978
rect 132038 154294 132094 154350
rect 132162 154294 132218 154350
rect 132038 154170 132094 154226
rect 132162 154170 132218 154226
rect 132038 154046 132094 154102
rect 132162 154046 132218 154102
rect 132038 153922 132094 153978
rect 132162 153922 132218 153978
rect 162758 154294 162814 154350
rect 162882 154294 162938 154350
rect 162758 154170 162814 154226
rect 162882 154170 162938 154226
rect 162758 154046 162814 154102
rect 162882 154046 162938 154102
rect 162758 153922 162814 153978
rect 162882 153922 162938 153978
rect 193478 154294 193534 154350
rect 193602 154294 193658 154350
rect 193478 154170 193534 154226
rect 193602 154170 193658 154226
rect 193478 154046 193534 154102
rect 193602 154046 193658 154102
rect 193478 153922 193534 153978
rect 193602 153922 193658 153978
rect 224198 154294 224254 154350
rect 224322 154294 224378 154350
rect 224198 154170 224254 154226
rect 224322 154170 224378 154226
rect 224198 154046 224254 154102
rect 224322 154046 224378 154102
rect 224198 153922 224254 153978
rect 224322 153922 224378 153978
rect 254918 154294 254974 154350
rect 255042 154294 255098 154350
rect 254918 154170 254974 154226
rect 255042 154170 255098 154226
rect 254918 154046 254974 154102
rect 255042 154046 255098 154102
rect 254918 153922 254974 153978
rect 255042 153922 255098 153978
rect 285638 154294 285694 154350
rect 285762 154294 285818 154350
rect 285638 154170 285694 154226
rect 285762 154170 285818 154226
rect 285638 154046 285694 154102
rect 285762 154046 285818 154102
rect 285638 153922 285694 153978
rect 285762 153922 285818 153978
rect 316358 154294 316414 154350
rect 316482 154294 316538 154350
rect 316358 154170 316414 154226
rect 316482 154170 316538 154226
rect 316358 154046 316414 154102
rect 316482 154046 316538 154102
rect 316358 153922 316414 153978
rect 316482 153922 316538 153978
rect 347078 154294 347134 154350
rect 347202 154294 347258 154350
rect 347078 154170 347134 154226
rect 347202 154170 347258 154226
rect 347078 154046 347134 154102
rect 347202 154046 347258 154102
rect 347078 153922 347134 153978
rect 347202 153922 347258 153978
rect 377798 154294 377854 154350
rect 377922 154294 377978 154350
rect 377798 154170 377854 154226
rect 377922 154170 377978 154226
rect 377798 154046 377854 154102
rect 377922 154046 377978 154102
rect 377798 153922 377854 153978
rect 377922 153922 377978 153978
rect 408518 154294 408574 154350
rect 408642 154294 408698 154350
rect 408518 154170 408574 154226
rect 408642 154170 408698 154226
rect 408518 154046 408574 154102
rect 408642 154046 408698 154102
rect 408518 153922 408574 153978
rect 408642 153922 408698 153978
rect 439238 154294 439294 154350
rect 439362 154294 439418 154350
rect 439238 154170 439294 154226
rect 439362 154170 439418 154226
rect 439238 154046 439294 154102
rect 439362 154046 439418 154102
rect 439238 153922 439294 153978
rect 439362 153922 439418 153978
rect 469958 154294 470014 154350
rect 470082 154294 470138 154350
rect 469958 154170 470014 154226
rect 470082 154170 470138 154226
rect 469958 154046 470014 154102
rect 470082 154046 470138 154102
rect 469958 153922 470014 153978
rect 470082 153922 470138 153978
rect 500678 154294 500734 154350
rect 500802 154294 500858 154350
rect 500678 154170 500734 154226
rect 500802 154170 500858 154226
rect 500678 154046 500734 154102
rect 500802 154046 500858 154102
rect 500678 153922 500734 153978
rect 500802 153922 500858 153978
rect 24518 148294 24574 148350
rect 24642 148294 24698 148350
rect 24518 148170 24574 148226
rect 24642 148170 24698 148226
rect 24518 148046 24574 148102
rect 24642 148046 24698 148102
rect 24518 147922 24574 147978
rect 24642 147922 24698 147978
rect 55238 148294 55294 148350
rect 55362 148294 55418 148350
rect 55238 148170 55294 148226
rect 55362 148170 55418 148226
rect 55238 148046 55294 148102
rect 55362 148046 55418 148102
rect 55238 147922 55294 147978
rect 55362 147922 55418 147978
rect 85958 148294 86014 148350
rect 86082 148294 86138 148350
rect 85958 148170 86014 148226
rect 86082 148170 86138 148226
rect 85958 148046 86014 148102
rect 86082 148046 86138 148102
rect 85958 147922 86014 147978
rect 86082 147922 86138 147978
rect 116678 148294 116734 148350
rect 116802 148294 116858 148350
rect 116678 148170 116734 148226
rect 116802 148170 116858 148226
rect 116678 148046 116734 148102
rect 116802 148046 116858 148102
rect 116678 147922 116734 147978
rect 116802 147922 116858 147978
rect 147398 148294 147454 148350
rect 147522 148294 147578 148350
rect 147398 148170 147454 148226
rect 147522 148170 147578 148226
rect 147398 148046 147454 148102
rect 147522 148046 147578 148102
rect 147398 147922 147454 147978
rect 147522 147922 147578 147978
rect 178118 148294 178174 148350
rect 178242 148294 178298 148350
rect 178118 148170 178174 148226
rect 178242 148170 178298 148226
rect 178118 148046 178174 148102
rect 178242 148046 178298 148102
rect 178118 147922 178174 147978
rect 178242 147922 178298 147978
rect 208838 148294 208894 148350
rect 208962 148294 209018 148350
rect 208838 148170 208894 148226
rect 208962 148170 209018 148226
rect 208838 148046 208894 148102
rect 208962 148046 209018 148102
rect 208838 147922 208894 147978
rect 208962 147922 209018 147978
rect 239558 148294 239614 148350
rect 239682 148294 239738 148350
rect 239558 148170 239614 148226
rect 239682 148170 239738 148226
rect 239558 148046 239614 148102
rect 239682 148046 239738 148102
rect 239558 147922 239614 147978
rect 239682 147922 239738 147978
rect 270278 148294 270334 148350
rect 270402 148294 270458 148350
rect 270278 148170 270334 148226
rect 270402 148170 270458 148226
rect 270278 148046 270334 148102
rect 270402 148046 270458 148102
rect 270278 147922 270334 147978
rect 270402 147922 270458 147978
rect 300998 148294 301054 148350
rect 301122 148294 301178 148350
rect 300998 148170 301054 148226
rect 301122 148170 301178 148226
rect 300998 148046 301054 148102
rect 301122 148046 301178 148102
rect 300998 147922 301054 147978
rect 301122 147922 301178 147978
rect 331718 148294 331774 148350
rect 331842 148294 331898 148350
rect 331718 148170 331774 148226
rect 331842 148170 331898 148226
rect 331718 148046 331774 148102
rect 331842 148046 331898 148102
rect 331718 147922 331774 147978
rect 331842 147922 331898 147978
rect 362438 148294 362494 148350
rect 362562 148294 362618 148350
rect 362438 148170 362494 148226
rect 362562 148170 362618 148226
rect 362438 148046 362494 148102
rect 362562 148046 362618 148102
rect 362438 147922 362494 147978
rect 362562 147922 362618 147978
rect 393158 148294 393214 148350
rect 393282 148294 393338 148350
rect 393158 148170 393214 148226
rect 393282 148170 393338 148226
rect 393158 148046 393214 148102
rect 393282 148046 393338 148102
rect 393158 147922 393214 147978
rect 393282 147922 393338 147978
rect 423878 148294 423934 148350
rect 424002 148294 424058 148350
rect 423878 148170 423934 148226
rect 424002 148170 424058 148226
rect 423878 148046 423934 148102
rect 424002 148046 424058 148102
rect 423878 147922 423934 147978
rect 424002 147922 424058 147978
rect 454598 148294 454654 148350
rect 454722 148294 454778 148350
rect 454598 148170 454654 148226
rect 454722 148170 454778 148226
rect 454598 148046 454654 148102
rect 454722 148046 454778 148102
rect 454598 147922 454654 147978
rect 454722 147922 454778 147978
rect 485318 148294 485374 148350
rect 485442 148294 485498 148350
rect 485318 148170 485374 148226
rect 485442 148170 485498 148226
rect 485318 148046 485374 148102
rect 485442 148046 485498 148102
rect 485318 147922 485374 147978
rect 485442 147922 485498 147978
rect 516038 148294 516094 148350
rect 516162 148294 516218 148350
rect 516038 148170 516094 148226
rect 516162 148170 516218 148226
rect 516038 148046 516094 148102
rect 516162 148046 516218 148102
rect 516038 147922 516094 147978
rect 516162 147922 516218 147978
rect 525250 148294 525306 148350
rect 525374 148294 525430 148350
rect 525498 148294 525554 148350
rect 525622 148294 525678 148350
rect 525250 148170 525306 148226
rect 525374 148170 525430 148226
rect 525498 148170 525554 148226
rect 525622 148170 525678 148226
rect 525250 148046 525306 148102
rect 525374 148046 525430 148102
rect 525498 148046 525554 148102
rect 525622 148046 525678 148102
rect 525250 147922 525306 147978
rect 525374 147922 525430 147978
rect 525498 147922 525554 147978
rect 525622 147922 525678 147978
rect 6970 136294 7026 136350
rect 7094 136294 7150 136350
rect 7218 136294 7274 136350
rect 7342 136294 7398 136350
rect 6970 136170 7026 136226
rect 7094 136170 7150 136226
rect 7218 136170 7274 136226
rect 7342 136170 7398 136226
rect 6970 136046 7026 136102
rect 7094 136046 7150 136102
rect 7218 136046 7274 136102
rect 7342 136046 7398 136102
rect 6970 135922 7026 135978
rect 7094 135922 7150 135978
rect 7218 135922 7274 135978
rect 7342 135922 7398 135978
rect 39878 136294 39934 136350
rect 40002 136294 40058 136350
rect 39878 136170 39934 136226
rect 40002 136170 40058 136226
rect 39878 136046 39934 136102
rect 40002 136046 40058 136102
rect 39878 135922 39934 135978
rect 40002 135922 40058 135978
rect 70598 136294 70654 136350
rect 70722 136294 70778 136350
rect 70598 136170 70654 136226
rect 70722 136170 70778 136226
rect 70598 136046 70654 136102
rect 70722 136046 70778 136102
rect 70598 135922 70654 135978
rect 70722 135922 70778 135978
rect 101318 136294 101374 136350
rect 101442 136294 101498 136350
rect 101318 136170 101374 136226
rect 101442 136170 101498 136226
rect 101318 136046 101374 136102
rect 101442 136046 101498 136102
rect 101318 135922 101374 135978
rect 101442 135922 101498 135978
rect 132038 136294 132094 136350
rect 132162 136294 132218 136350
rect 132038 136170 132094 136226
rect 132162 136170 132218 136226
rect 132038 136046 132094 136102
rect 132162 136046 132218 136102
rect 132038 135922 132094 135978
rect 132162 135922 132218 135978
rect 162758 136294 162814 136350
rect 162882 136294 162938 136350
rect 162758 136170 162814 136226
rect 162882 136170 162938 136226
rect 162758 136046 162814 136102
rect 162882 136046 162938 136102
rect 162758 135922 162814 135978
rect 162882 135922 162938 135978
rect 193478 136294 193534 136350
rect 193602 136294 193658 136350
rect 193478 136170 193534 136226
rect 193602 136170 193658 136226
rect 193478 136046 193534 136102
rect 193602 136046 193658 136102
rect 193478 135922 193534 135978
rect 193602 135922 193658 135978
rect 224198 136294 224254 136350
rect 224322 136294 224378 136350
rect 224198 136170 224254 136226
rect 224322 136170 224378 136226
rect 224198 136046 224254 136102
rect 224322 136046 224378 136102
rect 224198 135922 224254 135978
rect 224322 135922 224378 135978
rect 254918 136294 254974 136350
rect 255042 136294 255098 136350
rect 254918 136170 254974 136226
rect 255042 136170 255098 136226
rect 254918 136046 254974 136102
rect 255042 136046 255098 136102
rect 254918 135922 254974 135978
rect 255042 135922 255098 135978
rect 285638 136294 285694 136350
rect 285762 136294 285818 136350
rect 285638 136170 285694 136226
rect 285762 136170 285818 136226
rect 285638 136046 285694 136102
rect 285762 136046 285818 136102
rect 285638 135922 285694 135978
rect 285762 135922 285818 135978
rect 316358 136294 316414 136350
rect 316482 136294 316538 136350
rect 316358 136170 316414 136226
rect 316482 136170 316538 136226
rect 316358 136046 316414 136102
rect 316482 136046 316538 136102
rect 316358 135922 316414 135978
rect 316482 135922 316538 135978
rect 347078 136294 347134 136350
rect 347202 136294 347258 136350
rect 347078 136170 347134 136226
rect 347202 136170 347258 136226
rect 347078 136046 347134 136102
rect 347202 136046 347258 136102
rect 347078 135922 347134 135978
rect 347202 135922 347258 135978
rect 377798 136294 377854 136350
rect 377922 136294 377978 136350
rect 377798 136170 377854 136226
rect 377922 136170 377978 136226
rect 377798 136046 377854 136102
rect 377922 136046 377978 136102
rect 377798 135922 377854 135978
rect 377922 135922 377978 135978
rect 408518 136294 408574 136350
rect 408642 136294 408698 136350
rect 408518 136170 408574 136226
rect 408642 136170 408698 136226
rect 408518 136046 408574 136102
rect 408642 136046 408698 136102
rect 408518 135922 408574 135978
rect 408642 135922 408698 135978
rect 439238 136294 439294 136350
rect 439362 136294 439418 136350
rect 439238 136170 439294 136226
rect 439362 136170 439418 136226
rect 439238 136046 439294 136102
rect 439362 136046 439418 136102
rect 439238 135922 439294 135978
rect 439362 135922 439418 135978
rect 469958 136294 470014 136350
rect 470082 136294 470138 136350
rect 469958 136170 470014 136226
rect 470082 136170 470138 136226
rect 469958 136046 470014 136102
rect 470082 136046 470138 136102
rect 469958 135922 470014 135978
rect 470082 135922 470138 135978
rect 500678 136294 500734 136350
rect 500802 136294 500858 136350
rect 500678 136170 500734 136226
rect 500802 136170 500858 136226
rect 500678 136046 500734 136102
rect 500802 136046 500858 136102
rect 500678 135922 500734 135978
rect 500802 135922 500858 135978
rect 24518 130294 24574 130350
rect 24642 130294 24698 130350
rect 24518 130170 24574 130226
rect 24642 130170 24698 130226
rect 24518 130046 24574 130102
rect 24642 130046 24698 130102
rect 24518 129922 24574 129978
rect 24642 129922 24698 129978
rect 55238 130294 55294 130350
rect 55362 130294 55418 130350
rect 55238 130170 55294 130226
rect 55362 130170 55418 130226
rect 55238 130046 55294 130102
rect 55362 130046 55418 130102
rect 55238 129922 55294 129978
rect 55362 129922 55418 129978
rect 85958 130294 86014 130350
rect 86082 130294 86138 130350
rect 85958 130170 86014 130226
rect 86082 130170 86138 130226
rect 85958 130046 86014 130102
rect 86082 130046 86138 130102
rect 85958 129922 86014 129978
rect 86082 129922 86138 129978
rect 116678 130294 116734 130350
rect 116802 130294 116858 130350
rect 116678 130170 116734 130226
rect 116802 130170 116858 130226
rect 116678 130046 116734 130102
rect 116802 130046 116858 130102
rect 116678 129922 116734 129978
rect 116802 129922 116858 129978
rect 147398 130294 147454 130350
rect 147522 130294 147578 130350
rect 147398 130170 147454 130226
rect 147522 130170 147578 130226
rect 147398 130046 147454 130102
rect 147522 130046 147578 130102
rect 147398 129922 147454 129978
rect 147522 129922 147578 129978
rect 178118 130294 178174 130350
rect 178242 130294 178298 130350
rect 178118 130170 178174 130226
rect 178242 130170 178298 130226
rect 178118 130046 178174 130102
rect 178242 130046 178298 130102
rect 178118 129922 178174 129978
rect 178242 129922 178298 129978
rect 208838 130294 208894 130350
rect 208962 130294 209018 130350
rect 208838 130170 208894 130226
rect 208962 130170 209018 130226
rect 208838 130046 208894 130102
rect 208962 130046 209018 130102
rect 208838 129922 208894 129978
rect 208962 129922 209018 129978
rect 239558 130294 239614 130350
rect 239682 130294 239738 130350
rect 239558 130170 239614 130226
rect 239682 130170 239738 130226
rect 239558 130046 239614 130102
rect 239682 130046 239738 130102
rect 239558 129922 239614 129978
rect 239682 129922 239738 129978
rect 270278 130294 270334 130350
rect 270402 130294 270458 130350
rect 270278 130170 270334 130226
rect 270402 130170 270458 130226
rect 270278 130046 270334 130102
rect 270402 130046 270458 130102
rect 270278 129922 270334 129978
rect 270402 129922 270458 129978
rect 300998 130294 301054 130350
rect 301122 130294 301178 130350
rect 300998 130170 301054 130226
rect 301122 130170 301178 130226
rect 300998 130046 301054 130102
rect 301122 130046 301178 130102
rect 300998 129922 301054 129978
rect 301122 129922 301178 129978
rect 331718 130294 331774 130350
rect 331842 130294 331898 130350
rect 331718 130170 331774 130226
rect 331842 130170 331898 130226
rect 331718 130046 331774 130102
rect 331842 130046 331898 130102
rect 331718 129922 331774 129978
rect 331842 129922 331898 129978
rect 362438 130294 362494 130350
rect 362562 130294 362618 130350
rect 362438 130170 362494 130226
rect 362562 130170 362618 130226
rect 362438 130046 362494 130102
rect 362562 130046 362618 130102
rect 362438 129922 362494 129978
rect 362562 129922 362618 129978
rect 393158 130294 393214 130350
rect 393282 130294 393338 130350
rect 393158 130170 393214 130226
rect 393282 130170 393338 130226
rect 393158 130046 393214 130102
rect 393282 130046 393338 130102
rect 393158 129922 393214 129978
rect 393282 129922 393338 129978
rect 423878 130294 423934 130350
rect 424002 130294 424058 130350
rect 423878 130170 423934 130226
rect 424002 130170 424058 130226
rect 423878 130046 423934 130102
rect 424002 130046 424058 130102
rect 423878 129922 423934 129978
rect 424002 129922 424058 129978
rect 454598 130294 454654 130350
rect 454722 130294 454778 130350
rect 454598 130170 454654 130226
rect 454722 130170 454778 130226
rect 454598 130046 454654 130102
rect 454722 130046 454778 130102
rect 454598 129922 454654 129978
rect 454722 129922 454778 129978
rect 485318 130294 485374 130350
rect 485442 130294 485498 130350
rect 485318 130170 485374 130226
rect 485442 130170 485498 130226
rect 485318 130046 485374 130102
rect 485442 130046 485498 130102
rect 485318 129922 485374 129978
rect 485442 129922 485498 129978
rect 516038 130294 516094 130350
rect 516162 130294 516218 130350
rect 516038 130170 516094 130226
rect 516162 130170 516218 130226
rect 516038 130046 516094 130102
rect 516162 130046 516218 130102
rect 516038 129922 516094 129978
rect 516162 129922 516218 129978
rect 525250 130294 525306 130350
rect 525374 130294 525430 130350
rect 525498 130294 525554 130350
rect 525622 130294 525678 130350
rect 525250 130170 525306 130226
rect 525374 130170 525430 130226
rect 525498 130170 525554 130226
rect 525622 130170 525678 130226
rect 525250 130046 525306 130102
rect 525374 130046 525430 130102
rect 525498 130046 525554 130102
rect 525622 130046 525678 130102
rect 525250 129922 525306 129978
rect 525374 129922 525430 129978
rect 525498 129922 525554 129978
rect 525622 129922 525678 129978
rect 6970 118294 7026 118350
rect 7094 118294 7150 118350
rect 7218 118294 7274 118350
rect 7342 118294 7398 118350
rect 6970 118170 7026 118226
rect 7094 118170 7150 118226
rect 7218 118170 7274 118226
rect 7342 118170 7398 118226
rect 6970 118046 7026 118102
rect 7094 118046 7150 118102
rect 7218 118046 7274 118102
rect 7342 118046 7398 118102
rect 6970 117922 7026 117978
rect 7094 117922 7150 117978
rect 7218 117922 7274 117978
rect 7342 117922 7398 117978
rect 39878 118294 39934 118350
rect 40002 118294 40058 118350
rect 39878 118170 39934 118226
rect 40002 118170 40058 118226
rect 39878 118046 39934 118102
rect 40002 118046 40058 118102
rect 39878 117922 39934 117978
rect 40002 117922 40058 117978
rect 70598 118294 70654 118350
rect 70722 118294 70778 118350
rect 70598 118170 70654 118226
rect 70722 118170 70778 118226
rect 70598 118046 70654 118102
rect 70722 118046 70778 118102
rect 70598 117922 70654 117978
rect 70722 117922 70778 117978
rect 101318 118294 101374 118350
rect 101442 118294 101498 118350
rect 101318 118170 101374 118226
rect 101442 118170 101498 118226
rect 101318 118046 101374 118102
rect 101442 118046 101498 118102
rect 101318 117922 101374 117978
rect 101442 117922 101498 117978
rect 132038 118294 132094 118350
rect 132162 118294 132218 118350
rect 132038 118170 132094 118226
rect 132162 118170 132218 118226
rect 132038 118046 132094 118102
rect 132162 118046 132218 118102
rect 132038 117922 132094 117978
rect 132162 117922 132218 117978
rect 162758 118294 162814 118350
rect 162882 118294 162938 118350
rect 162758 118170 162814 118226
rect 162882 118170 162938 118226
rect 162758 118046 162814 118102
rect 162882 118046 162938 118102
rect 162758 117922 162814 117978
rect 162882 117922 162938 117978
rect 193478 118294 193534 118350
rect 193602 118294 193658 118350
rect 193478 118170 193534 118226
rect 193602 118170 193658 118226
rect 193478 118046 193534 118102
rect 193602 118046 193658 118102
rect 193478 117922 193534 117978
rect 193602 117922 193658 117978
rect 224198 118294 224254 118350
rect 224322 118294 224378 118350
rect 224198 118170 224254 118226
rect 224322 118170 224378 118226
rect 224198 118046 224254 118102
rect 224322 118046 224378 118102
rect 224198 117922 224254 117978
rect 224322 117922 224378 117978
rect 254918 118294 254974 118350
rect 255042 118294 255098 118350
rect 254918 118170 254974 118226
rect 255042 118170 255098 118226
rect 254918 118046 254974 118102
rect 255042 118046 255098 118102
rect 254918 117922 254974 117978
rect 255042 117922 255098 117978
rect 285638 118294 285694 118350
rect 285762 118294 285818 118350
rect 285638 118170 285694 118226
rect 285762 118170 285818 118226
rect 285638 118046 285694 118102
rect 285762 118046 285818 118102
rect 285638 117922 285694 117978
rect 285762 117922 285818 117978
rect 316358 118294 316414 118350
rect 316482 118294 316538 118350
rect 316358 118170 316414 118226
rect 316482 118170 316538 118226
rect 316358 118046 316414 118102
rect 316482 118046 316538 118102
rect 316358 117922 316414 117978
rect 316482 117922 316538 117978
rect 347078 118294 347134 118350
rect 347202 118294 347258 118350
rect 347078 118170 347134 118226
rect 347202 118170 347258 118226
rect 347078 118046 347134 118102
rect 347202 118046 347258 118102
rect 347078 117922 347134 117978
rect 347202 117922 347258 117978
rect 377798 118294 377854 118350
rect 377922 118294 377978 118350
rect 377798 118170 377854 118226
rect 377922 118170 377978 118226
rect 377798 118046 377854 118102
rect 377922 118046 377978 118102
rect 377798 117922 377854 117978
rect 377922 117922 377978 117978
rect 408518 118294 408574 118350
rect 408642 118294 408698 118350
rect 408518 118170 408574 118226
rect 408642 118170 408698 118226
rect 408518 118046 408574 118102
rect 408642 118046 408698 118102
rect 408518 117922 408574 117978
rect 408642 117922 408698 117978
rect 439238 118294 439294 118350
rect 439362 118294 439418 118350
rect 439238 118170 439294 118226
rect 439362 118170 439418 118226
rect 439238 118046 439294 118102
rect 439362 118046 439418 118102
rect 439238 117922 439294 117978
rect 439362 117922 439418 117978
rect 469958 118294 470014 118350
rect 470082 118294 470138 118350
rect 469958 118170 470014 118226
rect 470082 118170 470138 118226
rect 469958 118046 470014 118102
rect 470082 118046 470138 118102
rect 469958 117922 470014 117978
rect 470082 117922 470138 117978
rect 500678 118294 500734 118350
rect 500802 118294 500858 118350
rect 500678 118170 500734 118226
rect 500802 118170 500858 118226
rect 500678 118046 500734 118102
rect 500802 118046 500858 118102
rect 500678 117922 500734 117978
rect 500802 117922 500858 117978
rect 24518 112294 24574 112350
rect 24642 112294 24698 112350
rect 24518 112170 24574 112226
rect 24642 112170 24698 112226
rect 24518 112046 24574 112102
rect 24642 112046 24698 112102
rect 24518 111922 24574 111978
rect 24642 111922 24698 111978
rect 55238 112294 55294 112350
rect 55362 112294 55418 112350
rect 55238 112170 55294 112226
rect 55362 112170 55418 112226
rect 55238 112046 55294 112102
rect 55362 112046 55418 112102
rect 55238 111922 55294 111978
rect 55362 111922 55418 111978
rect 85958 112294 86014 112350
rect 86082 112294 86138 112350
rect 85958 112170 86014 112226
rect 86082 112170 86138 112226
rect 85958 112046 86014 112102
rect 86082 112046 86138 112102
rect 85958 111922 86014 111978
rect 86082 111922 86138 111978
rect 116678 112294 116734 112350
rect 116802 112294 116858 112350
rect 116678 112170 116734 112226
rect 116802 112170 116858 112226
rect 116678 112046 116734 112102
rect 116802 112046 116858 112102
rect 116678 111922 116734 111978
rect 116802 111922 116858 111978
rect 147398 112294 147454 112350
rect 147522 112294 147578 112350
rect 147398 112170 147454 112226
rect 147522 112170 147578 112226
rect 147398 112046 147454 112102
rect 147522 112046 147578 112102
rect 147398 111922 147454 111978
rect 147522 111922 147578 111978
rect 178118 112294 178174 112350
rect 178242 112294 178298 112350
rect 178118 112170 178174 112226
rect 178242 112170 178298 112226
rect 178118 112046 178174 112102
rect 178242 112046 178298 112102
rect 178118 111922 178174 111978
rect 178242 111922 178298 111978
rect 208838 112294 208894 112350
rect 208962 112294 209018 112350
rect 208838 112170 208894 112226
rect 208962 112170 209018 112226
rect 208838 112046 208894 112102
rect 208962 112046 209018 112102
rect 208838 111922 208894 111978
rect 208962 111922 209018 111978
rect 239558 112294 239614 112350
rect 239682 112294 239738 112350
rect 239558 112170 239614 112226
rect 239682 112170 239738 112226
rect 239558 112046 239614 112102
rect 239682 112046 239738 112102
rect 239558 111922 239614 111978
rect 239682 111922 239738 111978
rect 270278 112294 270334 112350
rect 270402 112294 270458 112350
rect 270278 112170 270334 112226
rect 270402 112170 270458 112226
rect 270278 112046 270334 112102
rect 270402 112046 270458 112102
rect 270278 111922 270334 111978
rect 270402 111922 270458 111978
rect 300998 112294 301054 112350
rect 301122 112294 301178 112350
rect 300998 112170 301054 112226
rect 301122 112170 301178 112226
rect 300998 112046 301054 112102
rect 301122 112046 301178 112102
rect 300998 111922 301054 111978
rect 301122 111922 301178 111978
rect 331718 112294 331774 112350
rect 331842 112294 331898 112350
rect 331718 112170 331774 112226
rect 331842 112170 331898 112226
rect 331718 112046 331774 112102
rect 331842 112046 331898 112102
rect 331718 111922 331774 111978
rect 331842 111922 331898 111978
rect 362438 112294 362494 112350
rect 362562 112294 362618 112350
rect 362438 112170 362494 112226
rect 362562 112170 362618 112226
rect 362438 112046 362494 112102
rect 362562 112046 362618 112102
rect 362438 111922 362494 111978
rect 362562 111922 362618 111978
rect 393158 112294 393214 112350
rect 393282 112294 393338 112350
rect 393158 112170 393214 112226
rect 393282 112170 393338 112226
rect 393158 112046 393214 112102
rect 393282 112046 393338 112102
rect 393158 111922 393214 111978
rect 393282 111922 393338 111978
rect 423878 112294 423934 112350
rect 424002 112294 424058 112350
rect 423878 112170 423934 112226
rect 424002 112170 424058 112226
rect 423878 112046 423934 112102
rect 424002 112046 424058 112102
rect 423878 111922 423934 111978
rect 424002 111922 424058 111978
rect 454598 112294 454654 112350
rect 454722 112294 454778 112350
rect 454598 112170 454654 112226
rect 454722 112170 454778 112226
rect 454598 112046 454654 112102
rect 454722 112046 454778 112102
rect 454598 111922 454654 111978
rect 454722 111922 454778 111978
rect 485318 112294 485374 112350
rect 485442 112294 485498 112350
rect 485318 112170 485374 112226
rect 485442 112170 485498 112226
rect 485318 112046 485374 112102
rect 485442 112046 485498 112102
rect 485318 111922 485374 111978
rect 485442 111922 485498 111978
rect 516038 112294 516094 112350
rect 516162 112294 516218 112350
rect 516038 112170 516094 112226
rect 516162 112170 516218 112226
rect 516038 112046 516094 112102
rect 516162 112046 516218 112102
rect 516038 111922 516094 111978
rect 516162 111922 516218 111978
rect 525250 112294 525306 112350
rect 525374 112294 525430 112350
rect 525498 112294 525554 112350
rect 525622 112294 525678 112350
rect 525250 112170 525306 112226
rect 525374 112170 525430 112226
rect 525498 112170 525554 112226
rect 525622 112170 525678 112226
rect 525250 112046 525306 112102
rect 525374 112046 525430 112102
rect 525498 112046 525554 112102
rect 525622 112046 525678 112102
rect 525250 111922 525306 111978
rect 525374 111922 525430 111978
rect 525498 111922 525554 111978
rect 525622 111922 525678 111978
rect 6970 100294 7026 100350
rect 7094 100294 7150 100350
rect 7218 100294 7274 100350
rect 7342 100294 7398 100350
rect 6970 100170 7026 100226
rect 7094 100170 7150 100226
rect 7218 100170 7274 100226
rect 7342 100170 7398 100226
rect 6970 100046 7026 100102
rect 7094 100046 7150 100102
rect 7218 100046 7274 100102
rect 7342 100046 7398 100102
rect 6970 99922 7026 99978
rect 7094 99922 7150 99978
rect 7218 99922 7274 99978
rect 7342 99922 7398 99978
rect 39878 100294 39934 100350
rect 40002 100294 40058 100350
rect 39878 100170 39934 100226
rect 40002 100170 40058 100226
rect 39878 100046 39934 100102
rect 40002 100046 40058 100102
rect 39878 99922 39934 99978
rect 40002 99922 40058 99978
rect 70598 100294 70654 100350
rect 70722 100294 70778 100350
rect 70598 100170 70654 100226
rect 70722 100170 70778 100226
rect 70598 100046 70654 100102
rect 70722 100046 70778 100102
rect 70598 99922 70654 99978
rect 70722 99922 70778 99978
rect 101318 100294 101374 100350
rect 101442 100294 101498 100350
rect 101318 100170 101374 100226
rect 101442 100170 101498 100226
rect 101318 100046 101374 100102
rect 101442 100046 101498 100102
rect 101318 99922 101374 99978
rect 101442 99922 101498 99978
rect 132038 100294 132094 100350
rect 132162 100294 132218 100350
rect 132038 100170 132094 100226
rect 132162 100170 132218 100226
rect 132038 100046 132094 100102
rect 132162 100046 132218 100102
rect 132038 99922 132094 99978
rect 132162 99922 132218 99978
rect 162758 100294 162814 100350
rect 162882 100294 162938 100350
rect 162758 100170 162814 100226
rect 162882 100170 162938 100226
rect 162758 100046 162814 100102
rect 162882 100046 162938 100102
rect 162758 99922 162814 99978
rect 162882 99922 162938 99978
rect 193478 100294 193534 100350
rect 193602 100294 193658 100350
rect 193478 100170 193534 100226
rect 193602 100170 193658 100226
rect 193478 100046 193534 100102
rect 193602 100046 193658 100102
rect 193478 99922 193534 99978
rect 193602 99922 193658 99978
rect 224198 100294 224254 100350
rect 224322 100294 224378 100350
rect 224198 100170 224254 100226
rect 224322 100170 224378 100226
rect 224198 100046 224254 100102
rect 224322 100046 224378 100102
rect 224198 99922 224254 99978
rect 224322 99922 224378 99978
rect 254918 100294 254974 100350
rect 255042 100294 255098 100350
rect 254918 100170 254974 100226
rect 255042 100170 255098 100226
rect 254918 100046 254974 100102
rect 255042 100046 255098 100102
rect 254918 99922 254974 99978
rect 255042 99922 255098 99978
rect 285638 100294 285694 100350
rect 285762 100294 285818 100350
rect 285638 100170 285694 100226
rect 285762 100170 285818 100226
rect 285638 100046 285694 100102
rect 285762 100046 285818 100102
rect 285638 99922 285694 99978
rect 285762 99922 285818 99978
rect 316358 100294 316414 100350
rect 316482 100294 316538 100350
rect 316358 100170 316414 100226
rect 316482 100170 316538 100226
rect 316358 100046 316414 100102
rect 316482 100046 316538 100102
rect 316358 99922 316414 99978
rect 316482 99922 316538 99978
rect 347078 100294 347134 100350
rect 347202 100294 347258 100350
rect 347078 100170 347134 100226
rect 347202 100170 347258 100226
rect 347078 100046 347134 100102
rect 347202 100046 347258 100102
rect 347078 99922 347134 99978
rect 347202 99922 347258 99978
rect 377798 100294 377854 100350
rect 377922 100294 377978 100350
rect 377798 100170 377854 100226
rect 377922 100170 377978 100226
rect 377798 100046 377854 100102
rect 377922 100046 377978 100102
rect 377798 99922 377854 99978
rect 377922 99922 377978 99978
rect 408518 100294 408574 100350
rect 408642 100294 408698 100350
rect 408518 100170 408574 100226
rect 408642 100170 408698 100226
rect 408518 100046 408574 100102
rect 408642 100046 408698 100102
rect 408518 99922 408574 99978
rect 408642 99922 408698 99978
rect 439238 100294 439294 100350
rect 439362 100294 439418 100350
rect 439238 100170 439294 100226
rect 439362 100170 439418 100226
rect 439238 100046 439294 100102
rect 439362 100046 439418 100102
rect 439238 99922 439294 99978
rect 439362 99922 439418 99978
rect 469958 100294 470014 100350
rect 470082 100294 470138 100350
rect 469958 100170 470014 100226
rect 470082 100170 470138 100226
rect 469958 100046 470014 100102
rect 470082 100046 470138 100102
rect 469958 99922 470014 99978
rect 470082 99922 470138 99978
rect 500678 100294 500734 100350
rect 500802 100294 500858 100350
rect 500678 100170 500734 100226
rect 500802 100170 500858 100226
rect 500678 100046 500734 100102
rect 500802 100046 500858 100102
rect 500678 99922 500734 99978
rect 500802 99922 500858 99978
rect 24518 94294 24574 94350
rect 24642 94294 24698 94350
rect 24518 94170 24574 94226
rect 24642 94170 24698 94226
rect 24518 94046 24574 94102
rect 24642 94046 24698 94102
rect 24518 93922 24574 93978
rect 24642 93922 24698 93978
rect 55238 94294 55294 94350
rect 55362 94294 55418 94350
rect 55238 94170 55294 94226
rect 55362 94170 55418 94226
rect 55238 94046 55294 94102
rect 55362 94046 55418 94102
rect 55238 93922 55294 93978
rect 55362 93922 55418 93978
rect 85958 94294 86014 94350
rect 86082 94294 86138 94350
rect 85958 94170 86014 94226
rect 86082 94170 86138 94226
rect 85958 94046 86014 94102
rect 86082 94046 86138 94102
rect 85958 93922 86014 93978
rect 86082 93922 86138 93978
rect 116678 94294 116734 94350
rect 116802 94294 116858 94350
rect 116678 94170 116734 94226
rect 116802 94170 116858 94226
rect 116678 94046 116734 94102
rect 116802 94046 116858 94102
rect 116678 93922 116734 93978
rect 116802 93922 116858 93978
rect 147398 94294 147454 94350
rect 147522 94294 147578 94350
rect 147398 94170 147454 94226
rect 147522 94170 147578 94226
rect 147398 94046 147454 94102
rect 147522 94046 147578 94102
rect 147398 93922 147454 93978
rect 147522 93922 147578 93978
rect 178118 94294 178174 94350
rect 178242 94294 178298 94350
rect 178118 94170 178174 94226
rect 178242 94170 178298 94226
rect 178118 94046 178174 94102
rect 178242 94046 178298 94102
rect 178118 93922 178174 93978
rect 178242 93922 178298 93978
rect 208838 94294 208894 94350
rect 208962 94294 209018 94350
rect 208838 94170 208894 94226
rect 208962 94170 209018 94226
rect 208838 94046 208894 94102
rect 208962 94046 209018 94102
rect 208838 93922 208894 93978
rect 208962 93922 209018 93978
rect 239558 94294 239614 94350
rect 239682 94294 239738 94350
rect 239558 94170 239614 94226
rect 239682 94170 239738 94226
rect 239558 94046 239614 94102
rect 239682 94046 239738 94102
rect 239558 93922 239614 93978
rect 239682 93922 239738 93978
rect 270278 94294 270334 94350
rect 270402 94294 270458 94350
rect 270278 94170 270334 94226
rect 270402 94170 270458 94226
rect 270278 94046 270334 94102
rect 270402 94046 270458 94102
rect 270278 93922 270334 93978
rect 270402 93922 270458 93978
rect 300998 94294 301054 94350
rect 301122 94294 301178 94350
rect 300998 94170 301054 94226
rect 301122 94170 301178 94226
rect 300998 94046 301054 94102
rect 301122 94046 301178 94102
rect 300998 93922 301054 93978
rect 301122 93922 301178 93978
rect 331718 94294 331774 94350
rect 331842 94294 331898 94350
rect 331718 94170 331774 94226
rect 331842 94170 331898 94226
rect 331718 94046 331774 94102
rect 331842 94046 331898 94102
rect 331718 93922 331774 93978
rect 331842 93922 331898 93978
rect 362438 94294 362494 94350
rect 362562 94294 362618 94350
rect 362438 94170 362494 94226
rect 362562 94170 362618 94226
rect 362438 94046 362494 94102
rect 362562 94046 362618 94102
rect 362438 93922 362494 93978
rect 362562 93922 362618 93978
rect 393158 94294 393214 94350
rect 393282 94294 393338 94350
rect 393158 94170 393214 94226
rect 393282 94170 393338 94226
rect 393158 94046 393214 94102
rect 393282 94046 393338 94102
rect 393158 93922 393214 93978
rect 393282 93922 393338 93978
rect 423878 94294 423934 94350
rect 424002 94294 424058 94350
rect 423878 94170 423934 94226
rect 424002 94170 424058 94226
rect 423878 94046 423934 94102
rect 424002 94046 424058 94102
rect 423878 93922 423934 93978
rect 424002 93922 424058 93978
rect 454598 94294 454654 94350
rect 454722 94294 454778 94350
rect 454598 94170 454654 94226
rect 454722 94170 454778 94226
rect 454598 94046 454654 94102
rect 454722 94046 454778 94102
rect 454598 93922 454654 93978
rect 454722 93922 454778 93978
rect 485318 94294 485374 94350
rect 485442 94294 485498 94350
rect 485318 94170 485374 94226
rect 485442 94170 485498 94226
rect 485318 94046 485374 94102
rect 485442 94046 485498 94102
rect 485318 93922 485374 93978
rect 485442 93922 485498 93978
rect 516038 94294 516094 94350
rect 516162 94294 516218 94350
rect 516038 94170 516094 94226
rect 516162 94170 516218 94226
rect 516038 94046 516094 94102
rect 516162 94046 516218 94102
rect 516038 93922 516094 93978
rect 516162 93922 516218 93978
rect 525250 94294 525306 94350
rect 525374 94294 525430 94350
rect 525498 94294 525554 94350
rect 525622 94294 525678 94350
rect 525250 94170 525306 94226
rect 525374 94170 525430 94226
rect 525498 94170 525554 94226
rect 525622 94170 525678 94226
rect 525250 94046 525306 94102
rect 525374 94046 525430 94102
rect 525498 94046 525554 94102
rect 525622 94046 525678 94102
rect 525250 93922 525306 93978
rect 525374 93922 525430 93978
rect 525498 93922 525554 93978
rect 525622 93922 525678 93978
rect 6970 82294 7026 82350
rect 7094 82294 7150 82350
rect 7218 82294 7274 82350
rect 7342 82294 7398 82350
rect 6970 82170 7026 82226
rect 7094 82170 7150 82226
rect 7218 82170 7274 82226
rect 7342 82170 7398 82226
rect 6970 82046 7026 82102
rect 7094 82046 7150 82102
rect 7218 82046 7274 82102
rect 7342 82046 7398 82102
rect 6970 81922 7026 81978
rect 7094 81922 7150 81978
rect 7218 81922 7274 81978
rect 7342 81922 7398 81978
rect 39878 82294 39934 82350
rect 40002 82294 40058 82350
rect 39878 82170 39934 82226
rect 40002 82170 40058 82226
rect 39878 82046 39934 82102
rect 40002 82046 40058 82102
rect 39878 81922 39934 81978
rect 40002 81922 40058 81978
rect 70598 82294 70654 82350
rect 70722 82294 70778 82350
rect 70598 82170 70654 82226
rect 70722 82170 70778 82226
rect 70598 82046 70654 82102
rect 70722 82046 70778 82102
rect 70598 81922 70654 81978
rect 70722 81922 70778 81978
rect 101318 82294 101374 82350
rect 101442 82294 101498 82350
rect 101318 82170 101374 82226
rect 101442 82170 101498 82226
rect 101318 82046 101374 82102
rect 101442 82046 101498 82102
rect 101318 81922 101374 81978
rect 101442 81922 101498 81978
rect 132038 82294 132094 82350
rect 132162 82294 132218 82350
rect 132038 82170 132094 82226
rect 132162 82170 132218 82226
rect 132038 82046 132094 82102
rect 132162 82046 132218 82102
rect 132038 81922 132094 81978
rect 132162 81922 132218 81978
rect 162758 82294 162814 82350
rect 162882 82294 162938 82350
rect 162758 82170 162814 82226
rect 162882 82170 162938 82226
rect 162758 82046 162814 82102
rect 162882 82046 162938 82102
rect 162758 81922 162814 81978
rect 162882 81922 162938 81978
rect 193478 82294 193534 82350
rect 193602 82294 193658 82350
rect 193478 82170 193534 82226
rect 193602 82170 193658 82226
rect 193478 82046 193534 82102
rect 193602 82046 193658 82102
rect 193478 81922 193534 81978
rect 193602 81922 193658 81978
rect 224198 82294 224254 82350
rect 224322 82294 224378 82350
rect 224198 82170 224254 82226
rect 224322 82170 224378 82226
rect 224198 82046 224254 82102
rect 224322 82046 224378 82102
rect 224198 81922 224254 81978
rect 224322 81922 224378 81978
rect 254918 82294 254974 82350
rect 255042 82294 255098 82350
rect 254918 82170 254974 82226
rect 255042 82170 255098 82226
rect 254918 82046 254974 82102
rect 255042 82046 255098 82102
rect 254918 81922 254974 81978
rect 255042 81922 255098 81978
rect 285638 82294 285694 82350
rect 285762 82294 285818 82350
rect 285638 82170 285694 82226
rect 285762 82170 285818 82226
rect 285638 82046 285694 82102
rect 285762 82046 285818 82102
rect 285638 81922 285694 81978
rect 285762 81922 285818 81978
rect 316358 82294 316414 82350
rect 316482 82294 316538 82350
rect 316358 82170 316414 82226
rect 316482 82170 316538 82226
rect 316358 82046 316414 82102
rect 316482 82046 316538 82102
rect 316358 81922 316414 81978
rect 316482 81922 316538 81978
rect 347078 82294 347134 82350
rect 347202 82294 347258 82350
rect 347078 82170 347134 82226
rect 347202 82170 347258 82226
rect 347078 82046 347134 82102
rect 347202 82046 347258 82102
rect 347078 81922 347134 81978
rect 347202 81922 347258 81978
rect 377798 82294 377854 82350
rect 377922 82294 377978 82350
rect 377798 82170 377854 82226
rect 377922 82170 377978 82226
rect 377798 82046 377854 82102
rect 377922 82046 377978 82102
rect 377798 81922 377854 81978
rect 377922 81922 377978 81978
rect 408518 82294 408574 82350
rect 408642 82294 408698 82350
rect 408518 82170 408574 82226
rect 408642 82170 408698 82226
rect 408518 82046 408574 82102
rect 408642 82046 408698 82102
rect 408518 81922 408574 81978
rect 408642 81922 408698 81978
rect 439238 82294 439294 82350
rect 439362 82294 439418 82350
rect 439238 82170 439294 82226
rect 439362 82170 439418 82226
rect 439238 82046 439294 82102
rect 439362 82046 439418 82102
rect 439238 81922 439294 81978
rect 439362 81922 439418 81978
rect 469958 82294 470014 82350
rect 470082 82294 470138 82350
rect 469958 82170 470014 82226
rect 470082 82170 470138 82226
rect 469958 82046 470014 82102
rect 470082 82046 470138 82102
rect 469958 81922 470014 81978
rect 470082 81922 470138 81978
rect 500678 82294 500734 82350
rect 500802 82294 500858 82350
rect 500678 82170 500734 82226
rect 500802 82170 500858 82226
rect 500678 82046 500734 82102
rect 500802 82046 500858 82102
rect 500678 81922 500734 81978
rect 500802 81922 500858 81978
rect 24518 76294 24574 76350
rect 24642 76294 24698 76350
rect 24518 76170 24574 76226
rect 24642 76170 24698 76226
rect 24518 76046 24574 76102
rect 24642 76046 24698 76102
rect 24518 75922 24574 75978
rect 24642 75922 24698 75978
rect 55238 76294 55294 76350
rect 55362 76294 55418 76350
rect 55238 76170 55294 76226
rect 55362 76170 55418 76226
rect 55238 76046 55294 76102
rect 55362 76046 55418 76102
rect 55238 75922 55294 75978
rect 55362 75922 55418 75978
rect 85958 76294 86014 76350
rect 86082 76294 86138 76350
rect 85958 76170 86014 76226
rect 86082 76170 86138 76226
rect 85958 76046 86014 76102
rect 86082 76046 86138 76102
rect 85958 75922 86014 75978
rect 86082 75922 86138 75978
rect 116678 76294 116734 76350
rect 116802 76294 116858 76350
rect 116678 76170 116734 76226
rect 116802 76170 116858 76226
rect 116678 76046 116734 76102
rect 116802 76046 116858 76102
rect 116678 75922 116734 75978
rect 116802 75922 116858 75978
rect 147398 76294 147454 76350
rect 147522 76294 147578 76350
rect 147398 76170 147454 76226
rect 147522 76170 147578 76226
rect 147398 76046 147454 76102
rect 147522 76046 147578 76102
rect 147398 75922 147454 75978
rect 147522 75922 147578 75978
rect 178118 76294 178174 76350
rect 178242 76294 178298 76350
rect 178118 76170 178174 76226
rect 178242 76170 178298 76226
rect 178118 76046 178174 76102
rect 178242 76046 178298 76102
rect 178118 75922 178174 75978
rect 178242 75922 178298 75978
rect 208838 76294 208894 76350
rect 208962 76294 209018 76350
rect 208838 76170 208894 76226
rect 208962 76170 209018 76226
rect 208838 76046 208894 76102
rect 208962 76046 209018 76102
rect 208838 75922 208894 75978
rect 208962 75922 209018 75978
rect 239558 76294 239614 76350
rect 239682 76294 239738 76350
rect 239558 76170 239614 76226
rect 239682 76170 239738 76226
rect 239558 76046 239614 76102
rect 239682 76046 239738 76102
rect 239558 75922 239614 75978
rect 239682 75922 239738 75978
rect 270278 76294 270334 76350
rect 270402 76294 270458 76350
rect 270278 76170 270334 76226
rect 270402 76170 270458 76226
rect 270278 76046 270334 76102
rect 270402 76046 270458 76102
rect 270278 75922 270334 75978
rect 270402 75922 270458 75978
rect 300998 76294 301054 76350
rect 301122 76294 301178 76350
rect 300998 76170 301054 76226
rect 301122 76170 301178 76226
rect 300998 76046 301054 76102
rect 301122 76046 301178 76102
rect 300998 75922 301054 75978
rect 301122 75922 301178 75978
rect 331718 76294 331774 76350
rect 331842 76294 331898 76350
rect 331718 76170 331774 76226
rect 331842 76170 331898 76226
rect 331718 76046 331774 76102
rect 331842 76046 331898 76102
rect 331718 75922 331774 75978
rect 331842 75922 331898 75978
rect 362438 76294 362494 76350
rect 362562 76294 362618 76350
rect 362438 76170 362494 76226
rect 362562 76170 362618 76226
rect 362438 76046 362494 76102
rect 362562 76046 362618 76102
rect 362438 75922 362494 75978
rect 362562 75922 362618 75978
rect 393158 76294 393214 76350
rect 393282 76294 393338 76350
rect 393158 76170 393214 76226
rect 393282 76170 393338 76226
rect 393158 76046 393214 76102
rect 393282 76046 393338 76102
rect 393158 75922 393214 75978
rect 393282 75922 393338 75978
rect 423878 76294 423934 76350
rect 424002 76294 424058 76350
rect 423878 76170 423934 76226
rect 424002 76170 424058 76226
rect 423878 76046 423934 76102
rect 424002 76046 424058 76102
rect 423878 75922 423934 75978
rect 424002 75922 424058 75978
rect 454598 76294 454654 76350
rect 454722 76294 454778 76350
rect 454598 76170 454654 76226
rect 454722 76170 454778 76226
rect 454598 76046 454654 76102
rect 454722 76046 454778 76102
rect 454598 75922 454654 75978
rect 454722 75922 454778 75978
rect 485318 76294 485374 76350
rect 485442 76294 485498 76350
rect 485318 76170 485374 76226
rect 485442 76170 485498 76226
rect 485318 76046 485374 76102
rect 485442 76046 485498 76102
rect 485318 75922 485374 75978
rect 485442 75922 485498 75978
rect 516038 76294 516094 76350
rect 516162 76294 516218 76350
rect 516038 76170 516094 76226
rect 516162 76170 516218 76226
rect 516038 76046 516094 76102
rect 516162 76046 516218 76102
rect 516038 75922 516094 75978
rect 516162 75922 516218 75978
rect 525250 76294 525306 76350
rect 525374 76294 525430 76350
rect 525498 76294 525554 76350
rect 525622 76294 525678 76350
rect 525250 76170 525306 76226
rect 525374 76170 525430 76226
rect 525498 76170 525554 76226
rect 525622 76170 525678 76226
rect 525250 76046 525306 76102
rect 525374 76046 525430 76102
rect 525498 76046 525554 76102
rect 525622 76046 525678 76102
rect 525250 75922 525306 75978
rect 525374 75922 525430 75978
rect 525498 75922 525554 75978
rect 525622 75922 525678 75978
rect 6970 64294 7026 64350
rect 7094 64294 7150 64350
rect 7218 64294 7274 64350
rect 7342 64294 7398 64350
rect 6970 64170 7026 64226
rect 7094 64170 7150 64226
rect 7218 64170 7274 64226
rect 7342 64170 7398 64226
rect 6970 64046 7026 64102
rect 7094 64046 7150 64102
rect 7218 64046 7274 64102
rect 7342 64046 7398 64102
rect 6970 63922 7026 63978
rect 7094 63922 7150 63978
rect 7218 63922 7274 63978
rect 7342 63922 7398 63978
rect 39878 64294 39934 64350
rect 40002 64294 40058 64350
rect 39878 64170 39934 64226
rect 40002 64170 40058 64226
rect 39878 64046 39934 64102
rect 40002 64046 40058 64102
rect 39878 63922 39934 63978
rect 40002 63922 40058 63978
rect 70598 64294 70654 64350
rect 70722 64294 70778 64350
rect 70598 64170 70654 64226
rect 70722 64170 70778 64226
rect 70598 64046 70654 64102
rect 70722 64046 70778 64102
rect 70598 63922 70654 63978
rect 70722 63922 70778 63978
rect 101318 64294 101374 64350
rect 101442 64294 101498 64350
rect 101318 64170 101374 64226
rect 101442 64170 101498 64226
rect 101318 64046 101374 64102
rect 101442 64046 101498 64102
rect 101318 63922 101374 63978
rect 101442 63922 101498 63978
rect 132038 64294 132094 64350
rect 132162 64294 132218 64350
rect 132038 64170 132094 64226
rect 132162 64170 132218 64226
rect 132038 64046 132094 64102
rect 132162 64046 132218 64102
rect 132038 63922 132094 63978
rect 132162 63922 132218 63978
rect 162758 64294 162814 64350
rect 162882 64294 162938 64350
rect 162758 64170 162814 64226
rect 162882 64170 162938 64226
rect 162758 64046 162814 64102
rect 162882 64046 162938 64102
rect 162758 63922 162814 63978
rect 162882 63922 162938 63978
rect 193478 64294 193534 64350
rect 193602 64294 193658 64350
rect 193478 64170 193534 64226
rect 193602 64170 193658 64226
rect 193478 64046 193534 64102
rect 193602 64046 193658 64102
rect 193478 63922 193534 63978
rect 193602 63922 193658 63978
rect 224198 64294 224254 64350
rect 224322 64294 224378 64350
rect 224198 64170 224254 64226
rect 224322 64170 224378 64226
rect 224198 64046 224254 64102
rect 224322 64046 224378 64102
rect 224198 63922 224254 63978
rect 224322 63922 224378 63978
rect 254918 64294 254974 64350
rect 255042 64294 255098 64350
rect 254918 64170 254974 64226
rect 255042 64170 255098 64226
rect 254918 64046 254974 64102
rect 255042 64046 255098 64102
rect 254918 63922 254974 63978
rect 255042 63922 255098 63978
rect 285638 64294 285694 64350
rect 285762 64294 285818 64350
rect 285638 64170 285694 64226
rect 285762 64170 285818 64226
rect 285638 64046 285694 64102
rect 285762 64046 285818 64102
rect 285638 63922 285694 63978
rect 285762 63922 285818 63978
rect 316358 64294 316414 64350
rect 316482 64294 316538 64350
rect 316358 64170 316414 64226
rect 316482 64170 316538 64226
rect 316358 64046 316414 64102
rect 316482 64046 316538 64102
rect 316358 63922 316414 63978
rect 316482 63922 316538 63978
rect 347078 64294 347134 64350
rect 347202 64294 347258 64350
rect 347078 64170 347134 64226
rect 347202 64170 347258 64226
rect 347078 64046 347134 64102
rect 347202 64046 347258 64102
rect 347078 63922 347134 63978
rect 347202 63922 347258 63978
rect 377798 64294 377854 64350
rect 377922 64294 377978 64350
rect 377798 64170 377854 64226
rect 377922 64170 377978 64226
rect 377798 64046 377854 64102
rect 377922 64046 377978 64102
rect 377798 63922 377854 63978
rect 377922 63922 377978 63978
rect 408518 64294 408574 64350
rect 408642 64294 408698 64350
rect 408518 64170 408574 64226
rect 408642 64170 408698 64226
rect 408518 64046 408574 64102
rect 408642 64046 408698 64102
rect 408518 63922 408574 63978
rect 408642 63922 408698 63978
rect 439238 64294 439294 64350
rect 439362 64294 439418 64350
rect 439238 64170 439294 64226
rect 439362 64170 439418 64226
rect 439238 64046 439294 64102
rect 439362 64046 439418 64102
rect 439238 63922 439294 63978
rect 439362 63922 439418 63978
rect 469958 64294 470014 64350
rect 470082 64294 470138 64350
rect 469958 64170 470014 64226
rect 470082 64170 470138 64226
rect 469958 64046 470014 64102
rect 470082 64046 470138 64102
rect 469958 63922 470014 63978
rect 470082 63922 470138 63978
rect 500678 64294 500734 64350
rect 500802 64294 500858 64350
rect 500678 64170 500734 64226
rect 500802 64170 500858 64226
rect 500678 64046 500734 64102
rect 500802 64046 500858 64102
rect 500678 63922 500734 63978
rect 500802 63922 500858 63978
rect 24518 58294 24574 58350
rect 24642 58294 24698 58350
rect 24518 58170 24574 58226
rect 24642 58170 24698 58226
rect 24518 58046 24574 58102
rect 24642 58046 24698 58102
rect 24518 57922 24574 57978
rect 24642 57922 24698 57978
rect 55238 58294 55294 58350
rect 55362 58294 55418 58350
rect 55238 58170 55294 58226
rect 55362 58170 55418 58226
rect 55238 58046 55294 58102
rect 55362 58046 55418 58102
rect 55238 57922 55294 57978
rect 55362 57922 55418 57978
rect 85958 58294 86014 58350
rect 86082 58294 86138 58350
rect 85958 58170 86014 58226
rect 86082 58170 86138 58226
rect 85958 58046 86014 58102
rect 86082 58046 86138 58102
rect 85958 57922 86014 57978
rect 86082 57922 86138 57978
rect 116678 58294 116734 58350
rect 116802 58294 116858 58350
rect 116678 58170 116734 58226
rect 116802 58170 116858 58226
rect 116678 58046 116734 58102
rect 116802 58046 116858 58102
rect 116678 57922 116734 57978
rect 116802 57922 116858 57978
rect 147398 58294 147454 58350
rect 147522 58294 147578 58350
rect 147398 58170 147454 58226
rect 147522 58170 147578 58226
rect 147398 58046 147454 58102
rect 147522 58046 147578 58102
rect 147398 57922 147454 57978
rect 147522 57922 147578 57978
rect 178118 58294 178174 58350
rect 178242 58294 178298 58350
rect 178118 58170 178174 58226
rect 178242 58170 178298 58226
rect 178118 58046 178174 58102
rect 178242 58046 178298 58102
rect 178118 57922 178174 57978
rect 178242 57922 178298 57978
rect 208838 58294 208894 58350
rect 208962 58294 209018 58350
rect 208838 58170 208894 58226
rect 208962 58170 209018 58226
rect 208838 58046 208894 58102
rect 208962 58046 209018 58102
rect 208838 57922 208894 57978
rect 208962 57922 209018 57978
rect 239558 58294 239614 58350
rect 239682 58294 239738 58350
rect 239558 58170 239614 58226
rect 239682 58170 239738 58226
rect 239558 58046 239614 58102
rect 239682 58046 239738 58102
rect 239558 57922 239614 57978
rect 239682 57922 239738 57978
rect 270278 58294 270334 58350
rect 270402 58294 270458 58350
rect 270278 58170 270334 58226
rect 270402 58170 270458 58226
rect 270278 58046 270334 58102
rect 270402 58046 270458 58102
rect 270278 57922 270334 57978
rect 270402 57922 270458 57978
rect 300998 58294 301054 58350
rect 301122 58294 301178 58350
rect 300998 58170 301054 58226
rect 301122 58170 301178 58226
rect 300998 58046 301054 58102
rect 301122 58046 301178 58102
rect 300998 57922 301054 57978
rect 301122 57922 301178 57978
rect 331718 58294 331774 58350
rect 331842 58294 331898 58350
rect 331718 58170 331774 58226
rect 331842 58170 331898 58226
rect 331718 58046 331774 58102
rect 331842 58046 331898 58102
rect 331718 57922 331774 57978
rect 331842 57922 331898 57978
rect 362438 58294 362494 58350
rect 362562 58294 362618 58350
rect 362438 58170 362494 58226
rect 362562 58170 362618 58226
rect 362438 58046 362494 58102
rect 362562 58046 362618 58102
rect 362438 57922 362494 57978
rect 362562 57922 362618 57978
rect 393158 58294 393214 58350
rect 393282 58294 393338 58350
rect 393158 58170 393214 58226
rect 393282 58170 393338 58226
rect 393158 58046 393214 58102
rect 393282 58046 393338 58102
rect 393158 57922 393214 57978
rect 393282 57922 393338 57978
rect 423878 58294 423934 58350
rect 424002 58294 424058 58350
rect 423878 58170 423934 58226
rect 424002 58170 424058 58226
rect 423878 58046 423934 58102
rect 424002 58046 424058 58102
rect 423878 57922 423934 57978
rect 424002 57922 424058 57978
rect 454598 58294 454654 58350
rect 454722 58294 454778 58350
rect 454598 58170 454654 58226
rect 454722 58170 454778 58226
rect 454598 58046 454654 58102
rect 454722 58046 454778 58102
rect 454598 57922 454654 57978
rect 454722 57922 454778 57978
rect 485318 58294 485374 58350
rect 485442 58294 485498 58350
rect 485318 58170 485374 58226
rect 485442 58170 485498 58226
rect 485318 58046 485374 58102
rect 485442 58046 485498 58102
rect 485318 57922 485374 57978
rect 485442 57922 485498 57978
rect 516038 58294 516094 58350
rect 516162 58294 516218 58350
rect 516038 58170 516094 58226
rect 516162 58170 516218 58226
rect 516038 58046 516094 58102
rect 516162 58046 516218 58102
rect 516038 57922 516094 57978
rect 516162 57922 516218 57978
rect 525250 58294 525306 58350
rect 525374 58294 525430 58350
rect 525498 58294 525554 58350
rect 525622 58294 525678 58350
rect 525250 58170 525306 58226
rect 525374 58170 525430 58226
rect 525498 58170 525554 58226
rect 525622 58170 525678 58226
rect 525250 58046 525306 58102
rect 525374 58046 525430 58102
rect 525498 58046 525554 58102
rect 525622 58046 525678 58102
rect 525250 57922 525306 57978
rect 525374 57922 525430 57978
rect 525498 57922 525554 57978
rect 525622 57922 525678 57978
rect 6970 46294 7026 46350
rect 7094 46294 7150 46350
rect 7218 46294 7274 46350
rect 7342 46294 7398 46350
rect 6970 46170 7026 46226
rect 7094 46170 7150 46226
rect 7218 46170 7274 46226
rect 7342 46170 7398 46226
rect 6970 46046 7026 46102
rect 7094 46046 7150 46102
rect 7218 46046 7274 46102
rect 7342 46046 7398 46102
rect 6970 45922 7026 45978
rect 7094 45922 7150 45978
rect 7218 45922 7274 45978
rect 7342 45922 7398 45978
rect 39878 46294 39934 46350
rect 40002 46294 40058 46350
rect 39878 46170 39934 46226
rect 40002 46170 40058 46226
rect 39878 46046 39934 46102
rect 40002 46046 40058 46102
rect 39878 45922 39934 45978
rect 40002 45922 40058 45978
rect 70598 46294 70654 46350
rect 70722 46294 70778 46350
rect 70598 46170 70654 46226
rect 70722 46170 70778 46226
rect 70598 46046 70654 46102
rect 70722 46046 70778 46102
rect 70598 45922 70654 45978
rect 70722 45922 70778 45978
rect 101318 46294 101374 46350
rect 101442 46294 101498 46350
rect 101318 46170 101374 46226
rect 101442 46170 101498 46226
rect 101318 46046 101374 46102
rect 101442 46046 101498 46102
rect 101318 45922 101374 45978
rect 101442 45922 101498 45978
rect 132038 46294 132094 46350
rect 132162 46294 132218 46350
rect 132038 46170 132094 46226
rect 132162 46170 132218 46226
rect 132038 46046 132094 46102
rect 132162 46046 132218 46102
rect 132038 45922 132094 45978
rect 132162 45922 132218 45978
rect 162758 46294 162814 46350
rect 162882 46294 162938 46350
rect 162758 46170 162814 46226
rect 162882 46170 162938 46226
rect 162758 46046 162814 46102
rect 162882 46046 162938 46102
rect 162758 45922 162814 45978
rect 162882 45922 162938 45978
rect 193478 46294 193534 46350
rect 193602 46294 193658 46350
rect 193478 46170 193534 46226
rect 193602 46170 193658 46226
rect 193478 46046 193534 46102
rect 193602 46046 193658 46102
rect 193478 45922 193534 45978
rect 193602 45922 193658 45978
rect 224198 46294 224254 46350
rect 224322 46294 224378 46350
rect 224198 46170 224254 46226
rect 224322 46170 224378 46226
rect 224198 46046 224254 46102
rect 224322 46046 224378 46102
rect 224198 45922 224254 45978
rect 224322 45922 224378 45978
rect 254918 46294 254974 46350
rect 255042 46294 255098 46350
rect 254918 46170 254974 46226
rect 255042 46170 255098 46226
rect 254918 46046 254974 46102
rect 255042 46046 255098 46102
rect 254918 45922 254974 45978
rect 255042 45922 255098 45978
rect 285638 46294 285694 46350
rect 285762 46294 285818 46350
rect 285638 46170 285694 46226
rect 285762 46170 285818 46226
rect 285638 46046 285694 46102
rect 285762 46046 285818 46102
rect 285638 45922 285694 45978
rect 285762 45922 285818 45978
rect 316358 46294 316414 46350
rect 316482 46294 316538 46350
rect 316358 46170 316414 46226
rect 316482 46170 316538 46226
rect 316358 46046 316414 46102
rect 316482 46046 316538 46102
rect 316358 45922 316414 45978
rect 316482 45922 316538 45978
rect 347078 46294 347134 46350
rect 347202 46294 347258 46350
rect 347078 46170 347134 46226
rect 347202 46170 347258 46226
rect 347078 46046 347134 46102
rect 347202 46046 347258 46102
rect 347078 45922 347134 45978
rect 347202 45922 347258 45978
rect 377798 46294 377854 46350
rect 377922 46294 377978 46350
rect 377798 46170 377854 46226
rect 377922 46170 377978 46226
rect 377798 46046 377854 46102
rect 377922 46046 377978 46102
rect 377798 45922 377854 45978
rect 377922 45922 377978 45978
rect 408518 46294 408574 46350
rect 408642 46294 408698 46350
rect 408518 46170 408574 46226
rect 408642 46170 408698 46226
rect 408518 46046 408574 46102
rect 408642 46046 408698 46102
rect 408518 45922 408574 45978
rect 408642 45922 408698 45978
rect 439238 46294 439294 46350
rect 439362 46294 439418 46350
rect 439238 46170 439294 46226
rect 439362 46170 439418 46226
rect 439238 46046 439294 46102
rect 439362 46046 439418 46102
rect 439238 45922 439294 45978
rect 439362 45922 439418 45978
rect 469958 46294 470014 46350
rect 470082 46294 470138 46350
rect 469958 46170 470014 46226
rect 470082 46170 470138 46226
rect 469958 46046 470014 46102
rect 470082 46046 470138 46102
rect 469958 45922 470014 45978
rect 470082 45922 470138 45978
rect 500678 46294 500734 46350
rect 500802 46294 500858 46350
rect 500678 46170 500734 46226
rect 500802 46170 500858 46226
rect 500678 46046 500734 46102
rect 500802 46046 500858 46102
rect 500678 45922 500734 45978
rect 500802 45922 500858 45978
rect 24518 40294 24574 40350
rect 24642 40294 24698 40350
rect 24518 40170 24574 40226
rect 24642 40170 24698 40226
rect 24518 40046 24574 40102
rect 24642 40046 24698 40102
rect 24518 39922 24574 39978
rect 24642 39922 24698 39978
rect 55238 40294 55294 40350
rect 55362 40294 55418 40350
rect 55238 40170 55294 40226
rect 55362 40170 55418 40226
rect 55238 40046 55294 40102
rect 55362 40046 55418 40102
rect 55238 39922 55294 39978
rect 55362 39922 55418 39978
rect 85958 40294 86014 40350
rect 86082 40294 86138 40350
rect 85958 40170 86014 40226
rect 86082 40170 86138 40226
rect 85958 40046 86014 40102
rect 86082 40046 86138 40102
rect 85958 39922 86014 39978
rect 86082 39922 86138 39978
rect 116678 40294 116734 40350
rect 116802 40294 116858 40350
rect 116678 40170 116734 40226
rect 116802 40170 116858 40226
rect 116678 40046 116734 40102
rect 116802 40046 116858 40102
rect 116678 39922 116734 39978
rect 116802 39922 116858 39978
rect 147398 40294 147454 40350
rect 147522 40294 147578 40350
rect 147398 40170 147454 40226
rect 147522 40170 147578 40226
rect 147398 40046 147454 40102
rect 147522 40046 147578 40102
rect 147398 39922 147454 39978
rect 147522 39922 147578 39978
rect 178118 40294 178174 40350
rect 178242 40294 178298 40350
rect 178118 40170 178174 40226
rect 178242 40170 178298 40226
rect 178118 40046 178174 40102
rect 178242 40046 178298 40102
rect 178118 39922 178174 39978
rect 178242 39922 178298 39978
rect 208838 40294 208894 40350
rect 208962 40294 209018 40350
rect 208838 40170 208894 40226
rect 208962 40170 209018 40226
rect 208838 40046 208894 40102
rect 208962 40046 209018 40102
rect 208838 39922 208894 39978
rect 208962 39922 209018 39978
rect 239558 40294 239614 40350
rect 239682 40294 239738 40350
rect 239558 40170 239614 40226
rect 239682 40170 239738 40226
rect 239558 40046 239614 40102
rect 239682 40046 239738 40102
rect 239558 39922 239614 39978
rect 239682 39922 239738 39978
rect 270278 40294 270334 40350
rect 270402 40294 270458 40350
rect 270278 40170 270334 40226
rect 270402 40170 270458 40226
rect 270278 40046 270334 40102
rect 270402 40046 270458 40102
rect 270278 39922 270334 39978
rect 270402 39922 270458 39978
rect 300998 40294 301054 40350
rect 301122 40294 301178 40350
rect 300998 40170 301054 40226
rect 301122 40170 301178 40226
rect 300998 40046 301054 40102
rect 301122 40046 301178 40102
rect 300998 39922 301054 39978
rect 301122 39922 301178 39978
rect 331718 40294 331774 40350
rect 331842 40294 331898 40350
rect 331718 40170 331774 40226
rect 331842 40170 331898 40226
rect 331718 40046 331774 40102
rect 331842 40046 331898 40102
rect 331718 39922 331774 39978
rect 331842 39922 331898 39978
rect 362438 40294 362494 40350
rect 362562 40294 362618 40350
rect 362438 40170 362494 40226
rect 362562 40170 362618 40226
rect 362438 40046 362494 40102
rect 362562 40046 362618 40102
rect 362438 39922 362494 39978
rect 362562 39922 362618 39978
rect 393158 40294 393214 40350
rect 393282 40294 393338 40350
rect 393158 40170 393214 40226
rect 393282 40170 393338 40226
rect 393158 40046 393214 40102
rect 393282 40046 393338 40102
rect 393158 39922 393214 39978
rect 393282 39922 393338 39978
rect 423878 40294 423934 40350
rect 424002 40294 424058 40350
rect 423878 40170 423934 40226
rect 424002 40170 424058 40226
rect 423878 40046 423934 40102
rect 424002 40046 424058 40102
rect 423878 39922 423934 39978
rect 424002 39922 424058 39978
rect 454598 40294 454654 40350
rect 454722 40294 454778 40350
rect 454598 40170 454654 40226
rect 454722 40170 454778 40226
rect 454598 40046 454654 40102
rect 454722 40046 454778 40102
rect 454598 39922 454654 39978
rect 454722 39922 454778 39978
rect 485318 40294 485374 40350
rect 485442 40294 485498 40350
rect 485318 40170 485374 40226
rect 485442 40170 485498 40226
rect 485318 40046 485374 40102
rect 485442 40046 485498 40102
rect 485318 39922 485374 39978
rect 485442 39922 485498 39978
rect 516038 40294 516094 40350
rect 516162 40294 516218 40350
rect 516038 40170 516094 40226
rect 516162 40170 516218 40226
rect 516038 40046 516094 40102
rect 516162 40046 516218 40102
rect 516038 39922 516094 39978
rect 516162 39922 516218 39978
rect 525250 40294 525306 40350
rect 525374 40294 525430 40350
rect 525498 40294 525554 40350
rect 525622 40294 525678 40350
rect 525250 40170 525306 40226
rect 525374 40170 525430 40226
rect 525498 40170 525554 40226
rect 525622 40170 525678 40226
rect 525250 40046 525306 40102
rect 525374 40046 525430 40102
rect 525498 40046 525554 40102
rect 525622 40046 525678 40102
rect 525250 39922 525306 39978
rect 525374 39922 525430 39978
rect 525498 39922 525554 39978
rect 525622 39922 525678 39978
rect 6970 28294 7026 28350
rect 7094 28294 7150 28350
rect 7218 28294 7274 28350
rect 7342 28294 7398 28350
rect 6970 28170 7026 28226
rect 7094 28170 7150 28226
rect 7218 28170 7274 28226
rect 7342 28170 7398 28226
rect 6970 28046 7026 28102
rect 7094 28046 7150 28102
rect 7218 28046 7274 28102
rect 7342 28046 7398 28102
rect 6970 27922 7026 27978
rect 7094 27922 7150 27978
rect 7218 27922 7274 27978
rect 7342 27922 7398 27978
rect 39878 28294 39934 28350
rect 40002 28294 40058 28350
rect 39878 28170 39934 28226
rect 40002 28170 40058 28226
rect 39878 28046 39934 28102
rect 40002 28046 40058 28102
rect 39878 27922 39934 27978
rect 40002 27922 40058 27978
rect 70598 28294 70654 28350
rect 70722 28294 70778 28350
rect 70598 28170 70654 28226
rect 70722 28170 70778 28226
rect 70598 28046 70654 28102
rect 70722 28046 70778 28102
rect 70598 27922 70654 27978
rect 70722 27922 70778 27978
rect 101318 28294 101374 28350
rect 101442 28294 101498 28350
rect 101318 28170 101374 28226
rect 101442 28170 101498 28226
rect 101318 28046 101374 28102
rect 101442 28046 101498 28102
rect 101318 27922 101374 27978
rect 101442 27922 101498 27978
rect 132038 28294 132094 28350
rect 132162 28294 132218 28350
rect 132038 28170 132094 28226
rect 132162 28170 132218 28226
rect 132038 28046 132094 28102
rect 132162 28046 132218 28102
rect 132038 27922 132094 27978
rect 132162 27922 132218 27978
rect 162758 28294 162814 28350
rect 162882 28294 162938 28350
rect 162758 28170 162814 28226
rect 162882 28170 162938 28226
rect 162758 28046 162814 28102
rect 162882 28046 162938 28102
rect 162758 27922 162814 27978
rect 162882 27922 162938 27978
rect 193478 28294 193534 28350
rect 193602 28294 193658 28350
rect 193478 28170 193534 28226
rect 193602 28170 193658 28226
rect 193478 28046 193534 28102
rect 193602 28046 193658 28102
rect 193478 27922 193534 27978
rect 193602 27922 193658 27978
rect 224198 28294 224254 28350
rect 224322 28294 224378 28350
rect 224198 28170 224254 28226
rect 224322 28170 224378 28226
rect 224198 28046 224254 28102
rect 224322 28046 224378 28102
rect 224198 27922 224254 27978
rect 224322 27922 224378 27978
rect 254918 28294 254974 28350
rect 255042 28294 255098 28350
rect 254918 28170 254974 28226
rect 255042 28170 255098 28226
rect 254918 28046 254974 28102
rect 255042 28046 255098 28102
rect 254918 27922 254974 27978
rect 255042 27922 255098 27978
rect 285638 28294 285694 28350
rect 285762 28294 285818 28350
rect 285638 28170 285694 28226
rect 285762 28170 285818 28226
rect 285638 28046 285694 28102
rect 285762 28046 285818 28102
rect 285638 27922 285694 27978
rect 285762 27922 285818 27978
rect 316358 28294 316414 28350
rect 316482 28294 316538 28350
rect 316358 28170 316414 28226
rect 316482 28170 316538 28226
rect 316358 28046 316414 28102
rect 316482 28046 316538 28102
rect 316358 27922 316414 27978
rect 316482 27922 316538 27978
rect 347078 28294 347134 28350
rect 347202 28294 347258 28350
rect 347078 28170 347134 28226
rect 347202 28170 347258 28226
rect 347078 28046 347134 28102
rect 347202 28046 347258 28102
rect 347078 27922 347134 27978
rect 347202 27922 347258 27978
rect 377798 28294 377854 28350
rect 377922 28294 377978 28350
rect 377798 28170 377854 28226
rect 377922 28170 377978 28226
rect 377798 28046 377854 28102
rect 377922 28046 377978 28102
rect 377798 27922 377854 27978
rect 377922 27922 377978 27978
rect 408518 28294 408574 28350
rect 408642 28294 408698 28350
rect 408518 28170 408574 28226
rect 408642 28170 408698 28226
rect 408518 28046 408574 28102
rect 408642 28046 408698 28102
rect 408518 27922 408574 27978
rect 408642 27922 408698 27978
rect 439238 28294 439294 28350
rect 439362 28294 439418 28350
rect 439238 28170 439294 28226
rect 439362 28170 439418 28226
rect 439238 28046 439294 28102
rect 439362 28046 439418 28102
rect 439238 27922 439294 27978
rect 439362 27922 439418 27978
rect 469958 28294 470014 28350
rect 470082 28294 470138 28350
rect 469958 28170 470014 28226
rect 470082 28170 470138 28226
rect 469958 28046 470014 28102
rect 470082 28046 470138 28102
rect 469958 27922 470014 27978
rect 470082 27922 470138 27978
rect 500678 28294 500734 28350
rect 500802 28294 500858 28350
rect 500678 28170 500734 28226
rect 500802 28170 500858 28226
rect 500678 28046 500734 28102
rect 500802 28046 500858 28102
rect 500678 27922 500734 27978
rect 500802 27922 500858 27978
rect 525250 22294 525306 22350
rect 525374 22294 525430 22350
rect 525498 22294 525554 22350
rect 525622 22294 525678 22350
rect 525250 22170 525306 22226
rect 525374 22170 525430 22226
rect 525498 22170 525554 22226
rect 525622 22170 525678 22226
rect 525250 22046 525306 22102
rect 525374 22046 525430 22102
rect 525498 22046 525554 22102
rect 525622 22046 525678 22102
rect 525250 21922 525306 21978
rect 525374 21922 525430 21978
rect 525498 21922 525554 21978
rect 525622 21922 525678 21978
rect 6970 10294 7026 10350
rect 7094 10294 7150 10350
rect 7218 10294 7274 10350
rect 7342 10294 7398 10350
rect 6970 10170 7026 10226
rect 7094 10170 7150 10226
rect 7218 10170 7274 10226
rect 7342 10170 7398 10226
rect 6970 10046 7026 10102
rect 7094 10046 7150 10102
rect 7218 10046 7274 10102
rect 7342 10046 7398 10102
rect 6970 9922 7026 9978
rect 7094 9922 7150 9978
rect 7218 9922 7274 9978
rect 7342 9922 7398 9978
rect 6970 -1176 7026 -1120
rect 7094 -1176 7150 -1120
rect 7218 -1176 7274 -1120
rect 7342 -1176 7398 -1120
rect 6970 -1300 7026 -1244
rect 7094 -1300 7150 -1244
rect 7218 -1300 7274 -1244
rect 7342 -1300 7398 -1244
rect 6970 -1424 7026 -1368
rect 7094 -1424 7150 -1368
rect 7218 -1424 7274 -1368
rect 7342 -1424 7398 -1368
rect 6970 -1548 7026 -1492
rect 7094 -1548 7150 -1492
rect 7218 -1548 7274 -1492
rect 7342 -1548 7398 -1492
rect 21250 4294 21306 4350
rect 21374 4294 21430 4350
rect 21498 4294 21554 4350
rect 21622 4294 21678 4350
rect 21250 4170 21306 4226
rect 21374 4170 21430 4226
rect 21498 4170 21554 4226
rect 21622 4170 21678 4226
rect 21250 4046 21306 4102
rect 21374 4046 21430 4102
rect 21498 4046 21554 4102
rect 21622 4046 21678 4102
rect 21250 3922 21306 3978
rect 21374 3922 21430 3978
rect 21498 3922 21554 3978
rect 21622 3922 21678 3978
rect 21250 -216 21306 -160
rect 21374 -216 21430 -160
rect 21498 -216 21554 -160
rect 21622 -216 21678 -160
rect 21250 -340 21306 -284
rect 21374 -340 21430 -284
rect 21498 -340 21554 -284
rect 21622 -340 21678 -284
rect 21250 -464 21306 -408
rect 21374 -464 21430 -408
rect 21498 -464 21554 -408
rect 21622 -464 21678 -408
rect 21250 -588 21306 -532
rect 21374 -588 21430 -532
rect 21498 -588 21554 -532
rect 21622 -588 21678 -532
rect 24970 10294 25026 10350
rect 25094 10294 25150 10350
rect 25218 10294 25274 10350
rect 25342 10294 25398 10350
rect 24970 10170 25026 10226
rect 25094 10170 25150 10226
rect 25218 10170 25274 10226
rect 25342 10170 25398 10226
rect 24970 10046 25026 10102
rect 25094 10046 25150 10102
rect 25218 10046 25274 10102
rect 25342 10046 25398 10102
rect 24970 9922 25026 9978
rect 25094 9922 25150 9978
rect 25218 9922 25274 9978
rect 25342 9922 25398 9978
rect 24970 -1176 25026 -1120
rect 25094 -1176 25150 -1120
rect 25218 -1176 25274 -1120
rect 25342 -1176 25398 -1120
rect 24970 -1300 25026 -1244
rect 25094 -1300 25150 -1244
rect 25218 -1300 25274 -1244
rect 25342 -1300 25398 -1244
rect 24970 -1424 25026 -1368
rect 25094 -1424 25150 -1368
rect 25218 -1424 25274 -1368
rect 25342 -1424 25398 -1368
rect 24970 -1548 25026 -1492
rect 25094 -1548 25150 -1492
rect 25218 -1548 25274 -1492
rect 25342 -1548 25398 -1492
rect 39250 4294 39306 4350
rect 39374 4294 39430 4350
rect 39498 4294 39554 4350
rect 39622 4294 39678 4350
rect 39250 4170 39306 4226
rect 39374 4170 39430 4226
rect 39498 4170 39554 4226
rect 39622 4170 39678 4226
rect 39250 4046 39306 4102
rect 39374 4046 39430 4102
rect 39498 4046 39554 4102
rect 39622 4046 39678 4102
rect 39250 3922 39306 3978
rect 39374 3922 39430 3978
rect 39498 3922 39554 3978
rect 39622 3922 39678 3978
rect 39250 -216 39306 -160
rect 39374 -216 39430 -160
rect 39498 -216 39554 -160
rect 39622 -216 39678 -160
rect 39250 -340 39306 -284
rect 39374 -340 39430 -284
rect 39498 -340 39554 -284
rect 39622 -340 39678 -284
rect 39250 -464 39306 -408
rect 39374 -464 39430 -408
rect 39498 -464 39554 -408
rect 39622 -464 39678 -408
rect 39250 -588 39306 -532
rect 39374 -588 39430 -532
rect 39498 -588 39554 -532
rect 39622 -588 39678 -532
rect 42970 10294 43026 10350
rect 43094 10294 43150 10350
rect 43218 10294 43274 10350
rect 43342 10294 43398 10350
rect 42970 10170 43026 10226
rect 43094 10170 43150 10226
rect 43218 10170 43274 10226
rect 43342 10170 43398 10226
rect 42970 10046 43026 10102
rect 43094 10046 43150 10102
rect 43218 10046 43274 10102
rect 43342 10046 43398 10102
rect 42970 9922 43026 9978
rect 43094 9922 43150 9978
rect 43218 9922 43274 9978
rect 43342 9922 43398 9978
rect 42970 -1176 43026 -1120
rect 43094 -1176 43150 -1120
rect 43218 -1176 43274 -1120
rect 43342 -1176 43398 -1120
rect 42970 -1300 43026 -1244
rect 43094 -1300 43150 -1244
rect 43218 -1300 43274 -1244
rect 43342 -1300 43398 -1244
rect 42970 -1424 43026 -1368
rect 43094 -1424 43150 -1368
rect 43218 -1424 43274 -1368
rect 43342 -1424 43398 -1368
rect 42970 -1548 43026 -1492
rect 43094 -1548 43150 -1492
rect 43218 -1548 43274 -1492
rect 43342 -1548 43398 -1492
rect 57250 4294 57306 4350
rect 57374 4294 57430 4350
rect 57498 4294 57554 4350
rect 57622 4294 57678 4350
rect 57250 4170 57306 4226
rect 57374 4170 57430 4226
rect 57498 4170 57554 4226
rect 57622 4170 57678 4226
rect 57250 4046 57306 4102
rect 57374 4046 57430 4102
rect 57498 4046 57554 4102
rect 57622 4046 57678 4102
rect 57250 3922 57306 3978
rect 57374 3922 57430 3978
rect 57498 3922 57554 3978
rect 57622 3922 57678 3978
rect 57250 -216 57306 -160
rect 57374 -216 57430 -160
rect 57498 -216 57554 -160
rect 57622 -216 57678 -160
rect 57250 -340 57306 -284
rect 57374 -340 57430 -284
rect 57498 -340 57554 -284
rect 57622 -340 57678 -284
rect 57250 -464 57306 -408
rect 57374 -464 57430 -408
rect 57498 -464 57554 -408
rect 57622 -464 57678 -408
rect 57250 -588 57306 -532
rect 57374 -588 57430 -532
rect 57498 -588 57554 -532
rect 57622 -588 57678 -532
rect 60970 10294 61026 10350
rect 61094 10294 61150 10350
rect 61218 10294 61274 10350
rect 61342 10294 61398 10350
rect 60970 10170 61026 10226
rect 61094 10170 61150 10226
rect 61218 10170 61274 10226
rect 61342 10170 61398 10226
rect 60970 10046 61026 10102
rect 61094 10046 61150 10102
rect 61218 10046 61274 10102
rect 61342 10046 61398 10102
rect 60970 9922 61026 9978
rect 61094 9922 61150 9978
rect 61218 9922 61274 9978
rect 61342 9922 61398 9978
rect 60970 -1176 61026 -1120
rect 61094 -1176 61150 -1120
rect 61218 -1176 61274 -1120
rect 61342 -1176 61398 -1120
rect 60970 -1300 61026 -1244
rect 61094 -1300 61150 -1244
rect 61218 -1300 61274 -1244
rect 61342 -1300 61398 -1244
rect 60970 -1424 61026 -1368
rect 61094 -1424 61150 -1368
rect 61218 -1424 61274 -1368
rect 61342 -1424 61398 -1368
rect 60970 -1548 61026 -1492
rect 61094 -1548 61150 -1492
rect 61218 -1548 61274 -1492
rect 61342 -1548 61398 -1492
rect 75250 4294 75306 4350
rect 75374 4294 75430 4350
rect 75498 4294 75554 4350
rect 75622 4294 75678 4350
rect 75250 4170 75306 4226
rect 75374 4170 75430 4226
rect 75498 4170 75554 4226
rect 75622 4170 75678 4226
rect 75250 4046 75306 4102
rect 75374 4046 75430 4102
rect 75498 4046 75554 4102
rect 75622 4046 75678 4102
rect 75250 3922 75306 3978
rect 75374 3922 75430 3978
rect 75498 3922 75554 3978
rect 75622 3922 75678 3978
rect 75250 -216 75306 -160
rect 75374 -216 75430 -160
rect 75498 -216 75554 -160
rect 75622 -216 75678 -160
rect 75250 -340 75306 -284
rect 75374 -340 75430 -284
rect 75498 -340 75554 -284
rect 75622 -340 75678 -284
rect 75250 -464 75306 -408
rect 75374 -464 75430 -408
rect 75498 -464 75554 -408
rect 75622 -464 75678 -408
rect 75250 -588 75306 -532
rect 75374 -588 75430 -532
rect 75498 -588 75554 -532
rect 75622 -588 75678 -532
rect 78970 10294 79026 10350
rect 79094 10294 79150 10350
rect 79218 10294 79274 10350
rect 79342 10294 79398 10350
rect 78970 10170 79026 10226
rect 79094 10170 79150 10226
rect 79218 10170 79274 10226
rect 79342 10170 79398 10226
rect 78970 10046 79026 10102
rect 79094 10046 79150 10102
rect 79218 10046 79274 10102
rect 79342 10046 79398 10102
rect 78970 9922 79026 9978
rect 79094 9922 79150 9978
rect 79218 9922 79274 9978
rect 79342 9922 79398 9978
rect 78970 -1176 79026 -1120
rect 79094 -1176 79150 -1120
rect 79218 -1176 79274 -1120
rect 79342 -1176 79398 -1120
rect 78970 -1300 79026 -1244
rect 79094 -1300 79150 -1244
rect 79218 -1300 79274 -1244
rect 79342 -1300 79398 -1244
rect 78970 -1424 79026 -1368
rect 79094 -1424 79150 -1368
rect 79218 -1424 79274 -1368
rect 79342 -1424 79398 -1368
rect 78970 -1548 79026 -1492
rect 79094 -1548 79150 -1492
rect 79218 -1548 79274 -1492
rect 79342 -1548 79398 -1492
rect 93250 4294 93306 4350
rect 93374 4294 93430 4350
rect 93498 4294 93554 4350
rect 93622 4294 93678 4350
rect 93250 4170 93306 4226
rect 93374 4170 93430 4226
rect 93498 4170 93554 4226
rect 93622 4170 93678 4226
rect 93250 4046 93306 4102
rect 93374 4046 93430 4102
rect 93498 4046 93554 4102
rect 93622 4046 93678 4102
rect 93250 3922 93306 3978
rect 93374 3922 93430 3978
rect 93498 3922 93554 3978
rect 93622 3922 93678 3978
rect 93250 -216 93306 -160
rect 93374 -216 93430 -160
rect 93498 -216 93554 -160
rect 93622 -216 93678 -160
rect 93250 -340 93306 -284
rect 93374 -340 93430 -284
rect 93498 -340 93554 -284
rect 93622 -340 93678 -284
rect 93250 -464 93306 -408
rect 93374 -464 93430 -408
rect 93498 -464 93554 -408
rect 93622 -464 93678 -408
rect 93250 -588 93306 -532
rect 93374 -588 93430 -532
rect 93498 -588 93554 -532
rect 93622 -588 93678 -532
rect 96970 10294 97026 10350
rect 97094 10294 97150 10350
rect 97218 10294 97274 10350
rect 97342 10294 97398 10350
rect 96970 10170 97026 10226
rect 97094 10170 97150 10226
rect 97218 10170 97274 10226
rect 97342 10170 97398 10226
rect 96970 10046 97026 10102
rect 97094 10046 97150 10102
rect 97218 10046 97274 10102
rect 97342 10046 97398 10102
rect 96970 9922 97026 9978
rect 97094 9922 97150 9978
rect 97218 9922 97274 9978
rect 97342 9922 97398 9978
rect 96970 -1176 97026 -1120
rect 97094 -1176 97150 -1120
rect 97218 -1176 97274 -1120
rect 97342 -1176 97398 -1120
rect 96970 -1300 97026 -1244
rect 97094 -1300 97150 -1244
rect 97218 -1300 97274 -1244
rect 97342 -1300 97398 -1244
rect 96970 -1424 97026 -1368
rect 97094 -1424 97150 -1368
rect 97218 -1424 97274 -1368
rect 97342 -1424 97398 -1368
rect 96970 -1548 97026 -1492
rect 97094 -1548 97150 -1492
rect 97218 -1548 97274 -1492
rect 97342 -1548 97398 -1492
rect 111250 4294 111306 4350
rect 111374 4294 111430 4350
rect 111498 4294 111554 4350
rect 111622 4294 111678 4350
rect 111250 4170 111306 4226
rect 111374 4170 111430 4226
rect 111498 4170 111554 4226
rect 111622 4170 111678 4226
rect 111250 4046 111306 4102
rect 111374 4046 111430 4102
rect 111498 4046 111554 4102
rect 111622 4046 111678 4102
rect 111250 3922 111306 3978
rect 111374 3922 111430 3978
rect 111498 3922 111554 3978
rect 111622 3922 111678 3978
rect 111250 -216 111306 -160
rect 111374 -216 111430 -160
rect 111498 -216 111554 -160
rect 111622 -216 111678 -160
rect 111250 -340 111306 -284
rect 111374 -340 111430 -284
rect 111498 -340 111554 -284
rect 111622 -340 111678 -284
rect 111250 -464 111306 -408
rect 111374 -464 111430 -408
rect 111498 -464 111554 -408
rect 111622 -464 111678 -408
rect 111250 -588 111306 -532
rect 111374 -588 111430 -532
rect 111498 -588 111554 -532
rect 111622 -588 111678 -532
rect 114970 10294 115026 10350
rect 115094 10294 115150 10350
rect 115218 10294 115274 10350
rect 115342 10294 115398 10350
rect 114970 10170 115026 10226
rect 115094 10170 115150 10226
rect 115218 10170 115274 10226
rect 115342 10170 115398 10226
rect 114970 10046 115026 10102
rect 115094 10046 115150 10102
rect 115218 10046 115274 10102
rect 115342 10046 115398 10102
rect 114970 9922 115026 9978
rect 115094 9922 115150 9978
rect 115218 9922 115274 9978
rect 115342 9922 115398 9978
rect 114970 -1176 115026 -1120
rect 115094 -1176 115150 -1120
rect 115218 -1176 115274 -1120
rect 115342 -1176 115398 -1120
rect 114970 -1300 115026 -1244
rect 115094 -1300 115150 -1244
rect 115218 -1300 115274 -1244
rect 115342 -1300 115398 -1244
rect 114970 -1424 115026 -1368
rect 115094 -1424 115150 -1368
rect 115218 -1424 115274 -1368
rect 115342 -1424 115398 -1368
rect 114970 -1548 115026 -1492
rect 115094 -1548 115150 -1492
rect 115218 -1548 115274 -1492
rect 115342 -1548 115398 -1492
rect 129250 4294 129306 4350
rect 129374 4294 129430 4350
rect 129498 4294 129554 4350
rect 129622 4294 129678 4350
rect 129250 4170 129306 4226
rect 129374 4170 129430 4226
rect 129498 4170 129554 4226
rect 129622 4170 129678 4226
rect 129250 4046 129306 4102
rect 129374 4046 129430 4102
rect 129498 4046 129554 4102
rect 129622 4046 129678 4102
rect 129250 3922 129306 3978
rect 129374 3922 129430 3978
rect 129498 3922 129554 3978
rect 129622 3922 129678 3978
rect 129250 -216 129306 -160
rect 129374 -216 129430 -160
rect 129498 -216 129554 -160
rect 129622 -216 129678 -160
rect 129250 -340 129306 -284
rect 129374 -340 129430 -284
rect 129498 -340 129554 -284
rect 129622 -340 129678 -284
rect 129250 -464 129306 -408
rect 129374 -464 129430 -408
rect 129498 -464 129554 -408
rect 129622 -464 129678 -408
rect 129250 -588 129306 -532
rect 129374 -588 129430 -532
rect 129498 -588 129554 -532
rect 129622 -588 129678 -532
rect 132970 10294 133026 10350
rect 133094 10294 133150 10350
rect 133218 10294 133274 10350
rect 133342 10294 133398 10350
rect 132970 10170 133026 10226
rect 133094 10170 133150 10226
rect 133218 10170 133274 10226
rect 133342 10170 133398 10226
rect 132970 10046 133026 10102
rect 133094 10046 133150 10102
rect 133218 10046 133274 10102
rect 133342 10046 133398 10102
rect 132970 9922 133026 9978
rect 133094 9922 133150 9978
rect 133218 9922 133274 9978
rect 133342 9922 133398 9978
rect 132970 -1176 133026 -1120
rect 133094 -1176 133150 -1120
rect 133218 -1176 133274 -1120
rect 133342 -1176 133398 -1120
rect 132970 -1300 133026 -1244
rect 133094 -1300 133150 -1244
rect 133218 -1300 133274 -1244
rect 133342 -1300 133398 -1244
rect 132970 -1424 133026 -1368
rect 133094 -1424 133150 -1368
rect 133218 -1424 133274 -1368
rect 133342 -1424 133398 -1368
rect 132970 -1548 133026 -1492
rect 133094 -1548 133150 -1492
rect 133218 -1548 133274 -1492
rect 133342 -1548 133398 -1492
rect 147250 4294 147306 4350
rect 147374 4294 147430 4350
rect 147498 4294 147554 4350
rect 147622 4294 147678 4350
rect 147250 4170 147306 4226
rect 147374 4170 147430 4226
rect 147498 4170 147554 4226
rect 147622 4170 147678 4226
rect 147250 4046 147306 4102
rect 147374 4046 147430 4102
rect 147498 4046 147554 4102
rect 147622 4046 147678 4102
rect 147250 3922 147306 3978
rect 147374 3922 147430 3978
rect 147498 3922 147554 3978
rect 147622 3922 147678 3978
rect 147250 -216 147306 -160
rect 147374 -216 147430 -160
rect 147498 -216 147554 -160
rect 147622 -216 147678 -160
rect 147250 -340 147306 -284
rect 147374 -340 147430 -284
rect 147498 -340 147554 -284
rect 147622 -340 147678 -284
rect 147250 -464 147306 -408
rect 147374 -464 147430 -408
rect 147498 -464 147554 -408
rect 147622 -464 147678 -408
rect 147250 -588 147306 -532
rect 147374 -588 147430 -532
rect 147498 -588 147554 -532
rect 147622 -588 147678 -532
rect 150970 10294 151026 10350
rect 151094 10294 151150 10350
rect 151218 10294 151274 10350
rect 151342 10294 151398 10350
rect 150970 10170 151026 10226
rect 151094 10170 151150 10226
rect 151218 10170 151274 10226
rect 151342 10170 151398 10226
rect 150970 10046 151026 10102
rect 151094 10046 151150 10102
rect 151218 10046 151274 10102
rect 151342 10046 151398 10102
rect 150970 9922 151026 9978
rect 151094 9922 151150 9978
rect 151218 9922 151274 9978
rect 151342 9922 151398 9978
rect 150970 -1176 151026 -1120
rect 151094 -1176 151150 -1120
rect 151218 -1176 151274 -1120
rect 151342 -1176 151398 -1120
rect 150970 -1300 151026 -1244
rect 151094 -1300 151150 -1244
rect 151218 -1300 151274 -1244
rect 151342 -1300 151398 -1244
rect 150970 -1424 151026 -1368
rect 151094 -1424 151150 -1368
rect 151218 -1424 151274 -1368
rect 151342 -1424 151398 -1368
rect 150970 -1548 151026 -1492
rect 151094 -1548 151150 -1492
rect 151218 -1548 151274 -1492
rect 151342 -1548 151398 -1492
rect 165250 4294 165306 4350
rect 165374 4294 165430 4350
rect 165498 4294 165554 4350
rect 165622 4294 165678 4350
rect 165250 4170 165306 4226
rect 165374 4170 165430 4226
rect 165498 4170 165554 4226
rect 165622 4170 165678 4226
rect 165250 4046 165306 4102
rect 165374 4046 165430 4102
rect 165498 4046 165554 4102
rect 165622 4046 165678 4102
rect 165250 3922 165306 3978
rect 165374 3922 165430 3978
rect 165498 3922 165554 3978
rect 165622 3922 165678 3978
rect 165250 -216 165306 -160
rect 165374 -216 165430 -160
rect 165498 -216 165554 -160
rect 165622 -216 165678 -160
rect 165250 -340 165306 -284
rect 165374 -340 165430 -284
rect 165498 -340 165554 -284
rect 165622 -340 165678 -284
rect 165250 -464 165306 -408
rect 165374 -464 165430 -408
rect 165498 -464 165554 -408
rect 165622 -464 165678 -408
rect 165250 -588 165306 -532
rect 165374 -588 165430 -532
rect 165498 -588 165554 -532
rect 165622 -588 165678 -532
rect 168970 10294 169026 10350
rect 169094 10294 169150 10350
rect 169218 10294 169274 10350
rect 169342 10294 169398 10350
rect 168970 10170 169026 10226
rect 169094 10170 169150 10226
rect 169218 10170 169274 10226
rect 169342 10170 169398 10226
rect 168970 10046 169026 10102
rect 169094 10046 169150 10102
rect 169218 10046 169274 10102
rect 169342 10046 169398 10102
rect 168970 9922 169026 9978
rect 169094 9922 169150 9978
rect 169218 9922 169274 9978
rect 169342 9922 169398 9978
rect 168970 -1176 169026 -1120
rect 169094 -1176 169150 -1120
rect 169218 -1176 169274 -1120
rect 169342 -1176 169398 -1120
rect 168970 -1300 169026 -1244
rect 169094 -1300 169150 -1244
rect 169218 -1300 169274 -1244
rect 169342 -1300 169398 -1244
rect 168970 -1424 169026 -1368
rect 169094 -1424 169150 -1368
rect 169218 -1424 169274 -1368
rect 169342 -1424 169398 -1368
rect 168970 -1548 169026 -1492
rect 169094 -1548 169150 -1492
rect 169218 -1548 169274 -1492
rect 169342 -1548 169398 -1492
rect 183250 4294 183306 4350
rect 183374 4294 183430 4350
rect 183498 4294 183554 4350
rect 183622 4294 183678 4350
rect 183250 4170 183306 4226
rect 183374 4170 183430 4226
rect 183498 4170 183554 4226
rect 183622 4170 183678 4226
rect 183250 4046 183306 4102
rect 183374 4046 183430 4102
rect 183498 4046 183554 4102
rect 183622 4046 183678 4102
rect 183250 3922 183306 3978
rect 183374 3922 183430 3978
rect 183498 3922 183554 3978
rect 183622 3922 183678 3978
rect 183250 -216 183306 -160
rect 183374 -216 183430 -160
rect 183498 -216 183554 -160
rect 183622 -216 183678 -160
rect 183250 -340 183306 -284
rect 183374 -340 183430 -284
rect 183498 -340 183554 -284
rect 183622 -340 183678 -284
rect 183250 -464 183306 -408
rect 183374 -464 183430 -408
rect 183498 -464 183554 -408
rect 183622 -464 183678 -408
rect 183250 -588 183306 -532
rect 183374 -588 183430 -532
rect 183498 -588 183554 -532
rect 183622 -588 183678 -532
rect 186970 10294 187026 10350
rect 187094 10294 187150 10350
rect 187218 10294 187274 10350
rect 187342 10294 187398 10350
rect 186970 10170 187026 10226
rect 187094 10170 187150 10226
rect 187218 10170 187274 10226
rect 187342 10170 187398 10226
rect 186970 10046 187026 10102
rect 187094 10046 187150 10102
rect 187218 10046 187274 10102
rect 187342 10046 187398 10102
rect 186970 9922 187026 9978
rect 187094 9922 187150 9978
rect 187218 9922 187274 9978
rect 187342 9922 187398 9978
rect 186970 -1176 187026 -1120
rect 187094 -1176 187150 -1120
rect 187218 -1176 187274 -1120
rect 187342 -1176 187398 -1120
rect 186970 -1300 187026 -1244
rect 187094 -1300 187150 -1244
rect 187218 -1300 187274 -1244
rect 187342 -1300 187398 -1244
rect 186970 -1424 187026 -1368
rect 187094 -1424 187150 -1368
rect 187218 -1424 187274 -1368
rect 187342 -1424 187398 -1368
rect 186970 -1548 187026 -1492
rect 187094 -1548 187150 -1492
rect 187218 -1548 187274 -1492
rect 187342 -1548 187398 -1492
rect 201250 4294 201306 4350
rect 201374 4294 201430 4350
rect 201498 4294 201554 4350
rect 201622 4294 201678 4350
rect 201250 4170 201306 4226
rect 201374 4170 201430 4226
rect 201498 4170 201554 4226
rect 201622 4170 201678 4226
rect 201250 4046 201306 4102
rect 201374 4046 201430 4102
rect 201498 4046 201554 4102
rect 201622 4046 201678 4102
rect 201250 3922 201306 3978
rect 201374 3922 201430 3978
rect 201498 3922 201554 3978
rect 201622 3922 201678 3978
rect 201250 -216 201306 -160
rect 201374 -216 201430 -160
rect 201498 -216 201554 -160
rect 201622 -216 201678 -160
rect 201250 -340 201306 -284
rect 201374 -340 201430 -284
rect 201498 -340 201554 -284
rect 201622 -340 201678 -284
rect 201250 -464 201306 -408
rect 201374 -464 201430 -408
rect 201498 -464 201554 -408
rect 201622 -464 201678 -408
rect 201250 -588 201306 -532
rect 201374 -588 201430 -532
rect 201498 -588 201554 -532
rect 201622 -588 201678 -532
rect 204970 10294 205026 10350
rect 205094 10294 205150 10350
rect 205218 10294 205274 10350
rect 205342 10294 205398 10350
rect 204970 10170 205026 10226
rect 205094 10170 205150 10226
rect 205218 10170 205274 10226
rect 205342 10170 205398 10226
rect 204970 10046 205026 10102
rect 205094 10046 205150 10102
rect 205218 10046 205274 10102
rect 205342 10046 205398 10102
rect 204970 9922 205026 9978
rect 205094 9922 205150 9978
rect 205218 9922 205274 9978
rect 205342 9922 205398 9978
rect 204970 -1176 205026 -1120
rect 205094 -1176 205150 -1120
rect 205218 -1176 205274 -1120
rect 205342 -1176 205398 -1120
rect 204970 -1300 205026 -1244
rect 205094 -1300 205150 -1244
rect 205218 -1300 205274 -1244
rect 205342 -1300 205398 -1244
rect 204970 -1424 205026 -1368
rect 205094 -1424 205150 -1368
rect 205218 -1424 205274 -1368
rect 205342 -1424 205398 -1368
rect 204970 -1548 205026 -1492
rect 205094 -1548 205150 -1492
rect 205218 -1548 205274 -1492
rect 205342 -1548 205398 -1492
rect 219250 4294 219306 4350
rect 219374 4294 219430 4350
rect 219498 4294 219554 4350
rect 219622 4294 219678 4350
rect 219250 4170 219306 4226
rect 219374 4170 219430 4226
rect 219498 4170 219554 4226
rect 219622 4170 219678 4226
rect 219250 4046 219306 4102
rect 219374 4046 219430 4102
rect 219498 4046 219554 4102
rect 219622 4046 219678 4102
rect 219250 3922 219306 3978
rect 219374 3922 219430 3978
rect 219498 3922 219554 3978
rect 219622 3922 219678 3978
rect 219250 -216 219306 -160
rect 219374 -216 219430 -160
rect 219498 -216 219554 -160
rect 219622 -216 219678 -160
rect 219250 -340 219306 -284
rect 219374 -340 219430 -284
rect 219498 -340 219554 -284
rect 219622 -340 219678 -284
rect 219250 -464 219306 -408
rect 219374 -464 219430 -408
rect 219498 -464 219554 -408
rect 219622 -464 219678 -408
rect 219250 -588 219306 -532
rect 219374 -588 219430 -532
rect 219498 -588 219554 -532
rect 219622 -588 219678 -532
rect 222970 10294 223026 10350
rect 223094 10294 223150 10350
rect 223218 10294 223274 10350
rect 223342 10294 223398 10350
rect 222970 10170 223026 10226
rect 223094 10170 223150 10226
rect 223218 10170 223274 10226
rect 223342 10170 223398 10226
rect 222970 10046 223026 10102
rect 223094 10046 223150 10102
rect 223218 10046 223274 10102
rect 223342 10046 223398 10102
rect 222970 9922 223026 9978
rect 223094 9922 223150 9978
rect 223218 9922 223274 9978
rect 223342 9922 223398 9978
rect 222970 -1176 223026 -1120
rect 223094 -1176 223150 -1120
rect 223218 -1176 223274 -1120
rect 223342 -1176 223398 -1120
rect 222970 -1300 223026 -1244
rect 223094 -1300 223150 -1244
rect 223218 -1300 223274 -1244
rect 223342 -1300 223398 -1244
rect 222970 -1424 223026 -1368
rect 223094 -1424 223150 -1368
rect 223218 -1424 223274 -1368
rect 223342 -1424 223398 -1368
rect 222970 -1548 223026 -1492
rect 223094 -1548 223150 -1492
rect 223218 -1548 223274 -1492
rect 223342 -1548 223398 -1492
rect 237250 4294 237306 4350
rect 237374 4294 237430 4350
rect 237498 4294 237554 4350
rect 237622 4294 237678 4350
rect 237250 4170 237306 4226
rect 237374 4170 237430 4226
rect 237498 4170 237554 4226
rect 237622 4170 237678 4226
rect 237250 4046 237306 4102
rect 237374 4046 237430 4102
rect 237498 4046 237554 4102
rect 237622 4046 237678 4102
rect 237250 3922 237306 3978
rect 237374 3922 237430 3978
rect 237498 3922 237554 3978
rect 237622 3922 237678 3978
rect 237250 -216 237306 -160
rect 237374 -216 237430 -160
rect 237498 -216 237554 -160
rect 237622 -216 237678 -160
rect 237250 -340 237306 -284
rect 237374 -340 237430 -284
rect 237498 -340 237554 -284
rect 237622 -340 237678 -284
rect 237250 -464 237306 -408
rect 237374 -464 237430 -408
rect 237498 -464 237554 -408
rect 237622 -464 237678 -408
rect 237250 -588 237306 -532
rect 237374 -588 237430 -532
rect 237498 -588 237554 -532
rect 237622 -588 237678 -532
rect 240970 10294 241026 10350
rect 241094 10294 241150 10350
rect 241218 10294 241274 10350
rect 241342 10294 241398 10350
rect 240970 10170 241026 10226
rect 241094 10170 241150 10226
rect 241218 10170 241274 10226
rect 241342 10170 241398 10226
rect 240970 10046 241026 10102
rect 241094 10046 241150 10102
rect 241218 10046 241274 10102
rect 241342 10046 241398 10102
rect 240970 9922 241026 9978
rect 241094 9922 241150 9978
rect 241218 9922 241274 9978
rect 241342 9922 241398 9978
rect 240970 -1176 241026 -1120
rect 241094 -1176 241150 -1120
rect 241218 -1176 241274 -1120
rect 241342 -1176 241398 -1120
rect 240970 -1300 241026 -1244
rect 241094 -1300 241150 -1244
rect 241218 -1300 241274 -1244
rect 241342 -1300 241398 -1244
rect 240970 -1424 241026 -1368
rect 241094 -1424 241150 -1368
rect 241218 -1424 241274 -1368
rect 241342 -1424 241398 -1368
rect 240970 -1548 241026 -1492
rect 241094 -1548 241150 -1492
rect 241218 -1548 241274 -1492
rect 241342 -1548 241398 -1492
rect 255250 4294 255306 4350
rect 255374 4294 255430 4350
rect 255498 4294 255554 4350
rect 255622 4294 255678 4350
rect 255250 4170 255306 4226
rect 255374 4170 255430 4226
rect 255498 4170 255554 4226
rect 255622 4170 255678 4226
rect 255250 4046 255306 4102
rect 255374 4046 255430 4102
rect 255498 4046 255554 4102
rect 255622 4046 255678 4102
rect 255250 3922 255306 3978
rect 255374 3922 255430 3978
rect 255498 3922 255554 3978
rect 255622 3922 255678 3978
rect 255250 -216 255306 -160
rect 255374 -216 255430 -160
rect 255498 -216 255554 -160
rect 255622 -216 255678 -160
rect 255250 -340 255306 -284
rect 255374 -340 255430 -284
rect 255498 -340 255554 -284
rect 255622 -340 255678 -284
rect 255250 -464 255306 -408
rect 255374 -464 255430 -408
rect 255498 -464 255554 -408
rect 255622 -464 255678 -408
rect 255250 -588 255306 -532
rect 255374 -588 255430 -532
rect 255498 -588 255554 -532
rect 255622 -588 255678 -532
rect 258970 10294 259026 10350
rect 259094 10294 259150 10350
rect 259218 10294 259274 10350
rect 259342 10294 259398 10350
rect 258970 10170 259026 10226
rect 259094 10170 259150 10226
rect 259218 10170 259274 10226
rect 259342 10170 259398 10226
rect 258970 10046 259026 10102
rect 259094 10046 259150 10102
rect 259218 10046 259274 10102
rect 259342 10046 259398 10102
rect 258970 9922 259026 9978
rect 259094 9922 259150 9978
rect 259218 9922 259274 9978
rect 259342 9922 259398 9978
rect 258970 -1176 259026 -1120
rect 259094 -1176 259150 -1120
rect 259218 -1176 259274 -1120
rect 259342 -1176 259398 -1120
rect 258970 -1300 259026 -1244
rect 259094 -1300 259150 -1244
rect 259218 -1300 259274 -1244
rect 259342 -1300 259398 -1244
rect 258970 -1424 259026 -1368
rect 259094 -1424 259150 -1368
rect 259218 -1424 259274 -1368
rect 259342 -1424 259398 -1368
rect 258970 -1548 259026 -1492
rect 259094 -1548 259150 -1492
rect 259218 -1548 259274 -1492
rect 259342 -1548 259398 -1492
rect 273250 4294 273306 4350
rect 273374 4294 273430 4350
rect 273498 4294 273554 4350
rect 273622 4294 273678 4350
rect 273250 4170 273306 4226
rect 273374 4170 273430 4226
rect 273498 4170 273554 4226
rect 273622 4170 273678 4226
rect 273250 4046 273306 4102
rect 273374 4046 273430 4102
rect 273498 4046 273554 4102
rect 273622 4046 273678 4102
rect 273250 3922 273306 3978
rect 273374 3922 273430 3978
rect 273498 3922 273554 3978
rect 273622 3922 273678 3978
rect 273250 -216 273306 -160
rect 273374 -216 273430 -160
rect 273498 -216 273554 -160
rect 273622 -216 273678 -160
rect 273250 -340 273306 -284
rect 273374 -340 273430 -284
rect 273498 -340 273554 -284
rect 273622 -340 273678 -284
rect 273250 -464 273306 -408
rect 273374 -464 273430 -408
rect 273498 -464 273554 -408
rect 273622 -464 273678 -408
rect 273250 -588 273306 -532
rect 273374 -588 273430 -532
rect 273498 -588 273554 -532
rect 273622 -588 273678 -532
rect 276970 10294 277026 10350
rect 277094 10294 277150 10350
rect 277218 10294 277274 10350
rect 277342 10294 277398 10350
rect 276970 10170 277026 10226
rect 277094 10170 277150 10226
rect 277218 10170 277274 10226
rect 277342 10170 277398 10226
rect 276970 10046 277026 10102
rect 277094 10046 277150 10102
rect 277218 10046 277274 10102
rect 277342 10046 277398 10102
rect 276970 9922 277026 9978
rect 277094 9922 277150 9978
rect 277218 9922 277274 9978
rect 277342 9922 277398 9978
rect 276970 -1176 277026 -1120
rect 277094 -1176 277150 -1120
rect 277218 -1176 277274 -1120
rect 277342 -1176 277398 -1120
rect 276970 -1300 277026 -1244
rect 277094 -1300 277150 -1244
rect 277218 -1300 277274 -1244
rect 277342 -1300 277398 -1244
rect 276970 -1424 277026 -1368
rect 277094 -1424 277150 -1368
rect 277218 -1424 277274 -1368
rect 277342 -1424 277398 -1368
rect 276970 -1548 277026 -1492
rect 277094 -1548 277150 -1492
rect 277218 -1548 277274 -1492
rect 277342 -1548 277398 -1492
rect 291250 4294 291306 4350
rect 291374 4294 291430 4350
rect 291498 4294 291554 4350
rect 291622 4294 291678 4350
rect 291250 4170 291306 4226
rect 291374 4170 291430 4226
rect 291498 4170 291554 4226
rect 291622 4170 291678 4226
rect 291250 4046 291306 4102
rect 291374 4046 291430 4102
rect 291498 4046 291554 4102
rect 291622 4046 291678 4102
rect 291250 3922 291306 3978
rect 291374 3922 291430 3978
rect 291498 3922 291554 3978
rect 291622 3922 291678 3978
rect 291250 -216 291306 -160
rect 291374 -216 291430 -160
rect 291498 -216 291554 -160
rect 291622 -216 291678 -160
rect 291250 -340 291306 -284
rect 291374 -340 291430 -284
rect 291498 -340 291554 -284
rect 291622 -340 291678 -284
rect 291250 -464 291306 -408
rect 291374 -464 291430 -408
rect 291498 -464 291554 -408
rect 291622 -464 291678 -408
rect 291250 -588 291306 -532
rect 291374 -588 291430 -532
rect 291498 -588 291554 -532
rect 291622 -588 291678 -532
rect 294970 10294 295026 10350
rect 295094 10294 295150 10350
rect 295218 10294 295274 10350
rect 295342 10294 295398 10350
rect 294970 10170 295026 10226
rect 295094 10170 295150 10226
rect 295218 10170 295274 10226
rect 295342 10170 295398 10226
rect 294970 10046 295026 10102
rect 295094 10046 295150 10102
rect 295218 10046 295274 10102
rect 295342 10046 295398 10102
rect 294970 9922 295026 9978
rect 295094 9922 295150 9978
rect 295218 9922 295274 9978
rect 295342 9922 295398 9978
rect 294970 -1176 295026 -1120
rect 295094 -1176 295150 -1120
rect 295218 -1176 295274 -1120
rect 295342 -1176 295398 -1120
rect 294970 -1300 295026 -1244
rect 295094 -1300 295150 -1244
rect 295218 -1300 295274 -1244
rect 295342 -1300 295398 -1244
rect 294970 -1424 295026 -1368
rect 295094 -1424 295150 -1368
rect 295218 -1424 295274 -1368
rect 295342 -1424 295398 -1368
rect 294970 -1548 295026 -1492
rect 295094 -1548 295150 -1492
rect 295218 -1548 295274 -1492
rect 295342 -1548 295398 -1492
rect 309250 4294 309306 4350
rect 309374 4294 309430 4350
rect 309498 4294 309554 4350
rect 309622 4294 309678 4350
rect 309250 4170 309306 4226
rect 309374 4170 309430 4226
rect 309498 4170 309554 4226
rect 309622 4170 309678 4226
rect 309250 4046 309306 4102
rect 309374 4046 309430 4102
rect 309498 4046 309554 4102
rect 309622 4046 309678 4102
rect 309250 3922 309306 3978
rect 309374 3922 309430 3978
rect 309498 3922 309554 3978
rect 309622 3922 309678 3978
rect 309250 -216 309306 -160
rect 309374 -216 309430 -160
rect 309498 -216 309554 -160
rect 309622 -216 309678 -160
rect 309250 -340 309306 -284
rect 309374 -340 309430 -284
rect 309498 -340 309554 -284
rect 309622 -340 309678 -284
rect 309250 -464 309306 -408
rect 309374 -464 309430 -408
rect 309498 -464 309554 -408
rect 309622 -464 309678 -408
rect 309250 -588 309306 -532
rect 309374 -588 309430 -532
rect 309498 -588 309554 -532
rect 309622 -588 309678 -532
rect 312970 10294 313026 10350
rect 313094 10294 313150 10350
rect 313218 10294 313274 10350
rect 313342 10294 313398 10350
rect 312970 10170 313026 10226
rect 313094 10170 313150 10226
rect 313218 10170 313274 10226
rect 313342 10170 313398 10226
rect 312970 10046 313026 10102
rect 313094 10046 313150 10102
rect 313218 10046 313274 10102
rect 313342 10046 313398 10102
rect 312970 9922 313026 9978
rect 313094 9922 313150 9978
rect 313218 9922 313274 9978
rect 313342 9922 313398 9978
rect 312970 -1176 313026 -1120
rect 313094 -1176 313150 -1120
rect 313218 -1176 313274 -1120
rect 313342 -1176 313398 -1120
rect 312970 -1300 313026 -1244
rect 313094 -1300 313150 -1244
rect 313218 -1300 313274 -1244
rect 313342 -1300 313398 -1244
rect 312970 -1424 313026 -1368
rect 313094 -1424 313150 -1368
rect 313218 -1424 313274 -1368
rect 313342 -1424 313398 -1368
rect 312970 -1548 313026 -1492
rect 313094 -1548 313150 -1492
rect 313218 -1548 313274 -1492
rect 313342 -1548 313398 -1492
rect 327250 4294 327306 4350
rect 327374 4294 327430 4350
rect 327498 4294 327554 4350
rect 327622 4294 327678 4350
rect 327250 4170 327306 4226
rect 327374 4170 327430 4226
rect 327498 4170 327554 4226
rect 327622 4170 327678 4226
rect 327250 4046 327306 4102
rect 327374 4046 327430 4102
rect 327498 4046 327554 4102
rect 327622 4046 327678 4102
rect 327250 3922 327306 3978
rect 327374 3922 327430 3978
rect 327498 3922 327554 3978
rect 327622 3922 327678 3978
rect 327250 -216 327306 -160
rect 327374 -216 327430 -160
rect 327498 -216 327554 -160
rect 327622 -216 327678 -160
rect 327250 -340 327306 -284
rect 327374 -340 327430 -284
rect 327498 -340 327554 -284
rect 327622 -340 327678 -284
rect 327250 -464 327306 -408
rect 327374 -464 327430 -408
rect 327498 -464 327554 -408
rect 327622 -464 327678 -408
rect 327250 -588 327306 -532
rect 327374 -588 327430 -532
rect 327498 -588 327554 -532
rect 327622 -588 327678 -532
rect 330970 10294 331026 10350
rect 331094 10294 331150 10350
rect 331218 10294 331274 10350
rect 331342 10294 331398 10350
rect 330970 10170 331026 10226
rect 331094 10170 331150 10226
rect 331218 10170 331274 10226
rect 331342 10170 331398 10226
rect 330970 10046 331026 10102
rect 331094 10046 331150 10102
rect 331218 10046 331274 10102
rect 331342 10046 331398 10102
rect 330970 9922 331026 9978
rect 331094 9922 331150 9978
rect 331218 9922 331274 9978
rect 331342 9922 331398 9978
rect 330970 -1176 331026 -1120
rect 331094 -1176 331150 -1120
rect 331218 -1176 331274 -1120
rect 331342 -1176 331398 -1120
rect 330970 -1300 331026 -1244
rect 331094 -1300 331150 -1244
rect 331218 -1300 331274 -1244
rect 331342 -1300 331398 -1244
rect 330970 -1424 331026 -1368
rect 331094 -1424 331150 -1368
rect 331218 -1424 331274 -1368
rect 331342 -1424 331398 -1368
rect 330970 -1548 331026 -1492
rect 331094 -1548 331150 -1492
rect 331218 -1548 331274 -1492
rect 331342 -1548 331398 -1492
rect 345250 4294 345306 4350
rect 345374 4294 345430 4350
rect 345498 4294 345554 4350
rect 345622 4294 345678 4350
rect 345250 4170 345306 4226
rect 345374 4170 345430 4226
rect 345498 4170 345554 4226
rect 345622 4170 345678 4226
rect 345250 4046 345306 4102
rect 345374 4046 345430 4102
rect 345498 4046 345554 4102
rect 345622 4046 345678 4102
rect 345250 3922 345306 3978
rect 345374 3922 345430 3978
rect 345498 3922 345554 3978
rect 345622 3922 345678 3978
rect 345250 -216 345306 -160
rect 345374 -216 345430 -160
rect 345498 -216 345554 -160
rect 345622 -216 345678 -160
rect 345250 -340 345306 -284
rect 345374 -340 345430 -284
rect 345498 -340 345554 -284
rect 345622 -340 345678 -284
rect 345250 -464 345306 -408
rect 345374 -464 345430 -408
rect 345498 -464 345554 -408
rect 345622 -464 345678 -408
rect 345250 -588 345306 -532
rect 345374 -588 345430 -532
rect 345498 -588 345554 -532
rect 345622 -588 345678 -532
rect 348970 10294 349026 10350
rect 349094 10294 349150 10350
rect 349218 10294 349274 10350
rect 349342 10294 349398 10350
rect 348970 10170 349026 10226
rect 349094 10170 349150 10226
rect 349218 10170 349274 10226
rect 349342 10170 349398 10226
rect 348970 10046 349026 10102
rect 349094 10046 349150 10102
rect 349218 10046 349274 10102
rect 349342 10046 349398 10102
rect 348970 9922 349026 9978
rect 349094 9922 349150 9978
rect 349218 9922 349274 9978
rect 349342 9922 349398 9978
rect 348970 -1176 349026 -1120
rect 349094 -1176 349150 -1120
rect 349218 -1176 349274 -1120
rect 349342 -1176 349398 -1120
rect 348970 -1300 349026 -1244
rect 349094 -1300 349150 -1244
rect 349218 -1300 349274 -1244
rect 349342 -1300 349398 -1244
rect 348970 -1424 349026 -1368
rect 349094 -1424 349150 -1368
rect 349218 -1424 349274 -1368
rect 349342 -1424 349398 -1368
rect 348970 -1548 349026 -1492
rect 349094 -1548 349150 -1492
rect 349218 -1548 349274 -1492
rect 349342 -1548 349398 -1492
rect 363250 4294 363306 4350
rect 363374 4294 363430 4350
rect 363498 4294 363554 4350
rect 363622 4294 363678 4350
rect 363250 4170 363306 4226
rect 363374 4170 363430 4226
rect 363498 4170 363554 4226
rect 363622 4170 363678 4226
rect 363250 4046 363306 4102
rect 363374 4046 363430 4102
rect 363498 4046 363554 4102
rect 363622 4046 363678 4102
rect 363250 3922 363306 3978
rect 363374 3922 363430 3978
rect 363498 3922 363554 3978
rect 363622 3922 363678 3978
rect 363250 -216 363306 -160
rect 363374 -216 363430 -160
rect 363498 -216 363554 -160
rect 363622 -216 363678 -160
rect 363250 -340 363306 -284
rect 363374 -340 363430 -284
rect 363498 -340 363554 -284
rect 363622 -340 363678 -284
rect 363250 -464 363306 -408
rect 363374 -464 363430 -408
rect 363498 -464 363554 -408
rect 363622 -464 363678 -408
rect 363250 -588 363306 -532
rect 363374 -588 363430 -532
rect 363498 -588 363554 -532
rect 363622 -588 363678 -532
rect 366970 10294 367026 10350
rect 367094 10294 367150 10350
rect 367218 10294 367274 10350
rect 367342 10294 367398 10350
rect 366970 10170 367026 10226
rect 367094 10170 367150 10226
rect 367218 10170 367274 10226
rect 367342 10170 367398 10226
rect 366970 10046 367026 10102
rect 367094 10046 367150 10102
rect 367218 10046 367274 10102
rect 367342 10046 367398 10102
rect 366970 9922 367026 9978
rect 367094 9922 367150 9978
rect 367218 9922 367274 9978
rect 367342 9922 367398 9978
rect 366970 -1176 367026 -1120
rect 367094 -1176 367150 -1120
rect 367218 -1176 367274 -1120
rect 367342 -1176 367398 -1120
rect 366970 -1300 367026 -1244
rect 367094 -1300 367150 -1244
rect 367218 -1300 367274 -1244
rect 367342 -1300 367398 -1244
rect 366970 -1424 367026 -1368
rect 367094 -1424 367150 -1368
rect 367218 -1424 367274 -1368
rect 367342 -1424 367398 -1368
rect 366970 -1548 367026 -1492
rect 367094 -1548 367150 -1492
rect 367218 -1548 367274 -1492
rect 367342 -1548 367398 -1492
rect 381250 4294 381306 4350
rect 381374 4294 381430 4350
rect 381498 4294 381554 4350
rect 381622 4294 381678 4350
rect 381250 4170 381306 4226
rect 381374 4170 381430 4226
rect 381498 4170 381554 4226
rect 381622 4170 381678 4226
rect 381250 4046 381306 4102
rect 381374 4046 381430 4102
rect 381498 4046 381554 4102
rect 381622 4046 381678 4102
rect 381250 3922 381306 3978
rect 381374 3922 381430 3978
rect 381498 3922 381554 3978
rect 381622 3922 381678 3978
rect 381250 -216 381306 -160
rect 381374 -216 381430 -160
rect 381498 -216 381554 -160
rect 381622 -216 381678 -160
rect 381250 -340 381306 -284
rect 381374 -340 381430 -284
rect 381498 -340 381554 -284
rect 381622 -340 381678 -284
rect 381250 -464 381306 -408
rect 381374 -464 381430 -408
rect 381498 -464 381554 -408
rect 381622 -464 381678 -408
rect 381250 -588 381306 -532
rect 381374 -588 381430 -532
rect 381498 -588 381554 -532
rect 381622 -588 381678 -532
rect 384970 10294 385026 10350
rect 385094 10294 385150 10350
rect 385218 10294 385274 10350
rect 385342 10294 385398 10350
rect 384970 10170 385026 10226
rect 385094 10170 385150 10226
rect 385218 10170 385274 10226
rect 385342 10170 385398 10226
rect 384970 10046 385026 10102
rect 385094 10046 385150 10102
rect 385218 10046 385274 10102
rect 385342 10046 385398 10102
rect 384970 9922 385026 9978
rect 385094 9922 385150 9978
rect 385218 9922 385274 9978
rect 385342 9922 385398 9978
rect 384970 -1176 385026 -1120
rect 385094 -1176 385150 -1120
rect 385218 -1176 385274 -1120
rect 385342 -1176 385398 -1120
rect 384970 -1300 385026 -1244
rect 385094 -1300 385150 -1244
rect 385218 -1300 385274 -1244
rect 385342 -1300 385398 -1244
rect 384970 -1424 385026 -1368
rect 385094 -1424 385150 -1368
rect 385218 -1424 385274 -1368
rect 385342 -1424 385398 -1368
rect 384970 -1548 385026 -1492
rect 385094 -1548 385150 -1492
rect 385218 -1548 385274 -1492
rect 385342 -1548 385398 -1492
rect 399250 4294 399306 4350
rect 399374 4294 399430 4350
rect 399498 4294 399554 4350
rect 399622 4294 399678 4350
rect 399250 4170 399306 4226
rect 399374 4170 399430 4226
rect 399498 4170 399554 4226
rect 399622 4170 399678 4226
rect 399250 4046 399306 4102
rect 399374 4046 399430 4102
rect 399498 4046 399554 4102
rect 399622 4046 399678 4102
rect 399250 3922 399306 3978
rect 399374 3922 399430 3978
rect 399498 3922 399554 3978
rect 399622 3922 399678 3978
rect 399250 -216 399306 -160
rect 399374 -216 399430 -160
rect 399498 -216 399554 -160
rect 399622 -216 399678 -160
rect 399250 -340 399306 -284
rect 399374 -340 399430 -284
rect 399498 -340 399554 -284
rect 399622 -340 399678 -284
rect 399250 -464 399306 -408
rect 399374 -464 399430 -408
rect 399498 -464 399554 -408
rect 399622 -464 399678 -408
rect 399250 -588 399306 -532
rect 399374 -588 399430 -532
rect 399498 -588 399554 -532
rect 399622 -588 399678 -532
rect 402970 10294 403026 10350
rect 403094 10294 403150 10350
rect 403218 10294 403274 10350
rect 403342 10294 403398 10350
rect 402970 10170 403026 10226
rect 403094 10170 403150 10226
rect 403218 10170 403274 10226
rect 403342 10170 403398 10226
rect 402970 10046 403026 10102
rect 403094 10046 403150 10102
rect 403218 10046 403274 10102
rect 403342 10046 403398 10102
rect 402970 9922 403026 9978
rect 403094 9922 403150 9978
rect 403218 9922 403274 9978
rect 403342 9922 403398 9978
rect 402970 -1176 403026 -1120
rect 403094 -1176 403150 -1120
rect 403218 -1176 403274 -1120
rect 403342 -1176 403398 -1120
rect 402970 -1300 403026 -1244
rect 403094 -1300 403150 -1244
rect 403218 -1300 403274 -1244
rect 403342 -1300 403398 -1244
rect 402970 -1424 403026 -1368
rect 403094 -1424 403150 -1368
rect 403218 -1424 403274 -1368
rect 403342 -1424 403398 -1368
rect 402970 -1548 403026 -1492
rect 403094 -1548 403150 -1492
rect 403218 -1548 403274 -1492
rect 403342 -1548 403398 -1492
rect 417250 4294 417306 4350
rect 417374 4294 417430 4350
rect 417498 4294 417554 4350
rect 417622 4294 417678 4350
rect 417250 4170 417306 4226
rect 417374 4170 417430 4226
rect 417498 4170 417554 4226
rect 417622 4170 417678 4226
rect 417250 4046 417306 4102
rect 417374 4046 417430 4102
rect 417498 4046 417554 4102
rect 417622 4046 417678 4102
rect 417250 3922 417306 3978
rect 417374 3922 417430 3978
rect 417498 3922 417554 3978
rect 417622 3922 417678 3978
rect 417250 -216 417306 -160
rect 417374 -216 417430 -160
rect 417498 -216 417554 -160
rect 417622 -216 417678 -160
rect 417250 -340 417306 -284
rect 417374 -340 417430 -284
rect 417498 -340 417554 -284
rect 417622 -340 417678 -284
rect 417250 -464 417306 -408
rect 417374 -464 417430 -408
rect 417498 -464 417554 -408
rect 417622 -464 417678 -408
rect 417250 -588 417306 -532
rect 417374 -588 417430 -532
rect 417498 -588 417554 -532
rect 417622 -588 417678 -532
rect 420970 10294 421026 10350
rect 421094 10294 421150 10350
rect 421218 10294 421274 10350
rect 421342 10294 421398 10350
rect 420970 10170 421026 10226
rect 421094 10170 421150 10226
rect 421218 10170 421274 10226
rect 421342 10170 421398 10226
rect 420970 10046 421026 10102
rect 421094 10046 421150 10102
rect 421218 10046 421274 10102
rect 421342 10046 421398 10102
rect 420970 9922 421026 9978
rect 421094 9922 421150 9978
rect 421218 9922 421274 9978
rect 421342 9922 421398 9978
rect 420970 -1176 421026 -1120
rect 421094 -1176 421150 -1120
rect 421218 -1176 421274 -1120
rect 421342 -1176 421398 -1120
rect 420970 -1300 421026 -1244
rect 421094 -1300 421150 -1244
rect 421218 -1300 421274 -1244
rect 421342 -1300 421398 -1244
rect 420970 -1424 421026 -1368
rect 421094 -1424 421150 -1368
rect 421218 -1424 421274 -1368
rect 421342 -1424 421398 -1368
rect 420970 -1548 421026 -1492
rect 421094 -1548 421150 -1492
rect 421218 -1548 421274 -1492
rect 421342 -1548 421398 -1492
rect 435250 4294 435306 4350
rect 435374 4294 435430 4350
rect 435498 4294 435554 4350
rect 435622 4294 435678 4350
rect 435250 4170 435306 4226
rect 435374 4170 435430 4226
rect 435498 4170 435554 4226
rect 435622 4170 435678 4226
rect 435250 4046 435306 4102
rect 435374 4046 435430 4102
rect 435498 4046 435554 4102
rect 435622 4046 435678 4102
rect 435250 3922 435306 3978
rect 435374 3922 435430 3978
rect 435498 3922 435554 3978
rect 435622 3922 435678 3978
rect 435250 -216 435306 -160
rect 435374 -216 435430 -160
rect 435498 -216 435554 -160
rect 435622 -216 435678 -160
rect 435250 -340 435306 -284
rect 435374 -340 435430 -284
rect 435498 -340 435554 -284
rect 435622 -340 435678 -284
rect 435250 -464 435306 -408
rect 435374 -464 435430 -408
rect 435498 -464 435554 -408
rect 435622 -464 435678 -408
rect 435250 -588 435306 -532
rect 435374 -588 435430 -532
rect 435498 -588 435554 -532
rect 435622 -588 435678 -532
rect 438970 10294 439026 10350
rect 439094 10294 439150 10350
rect 439218 10294 439274 10350
rect 439342 10294 439398 10350
rect 438970 10170 439026 10226
rect 439094 10170 439150 10226
rect 439218 10170 439274 10226
rect 439342 10170 439398 10226
rect 438970 10046 439026 10102
rect 439094 10046 439150 10102
rect 439218 10046 439274 10102
rect 439342 10046 439398 10102
rect 438970 9922 439026 9978
rect 439094 9922 439150 9978
rect 439218 9922 439274 9978
rect 439342 9922 439398 9978
rect 438970 -1176 439026 -1120
rect 439094 -1176 439150 -1120
rect 439218 -1176 439274 -1120
rect 439342 -1176 439398 -1120
rect 438970 -1300 439026 -1244
rect 439094 -1300 439150 -1244
rect 439218 -1300 439274 -1244
rect 439342 -1300 439398 -1244
rect 438970 -1424 439026 -1368
rect 439094 -1424 439150 -1368
rect 439218 -1424 439274 -1368
rect 439342 -1424 439398 -1368
rect 438970 -1548 439026 -1492
rect 439094 -1548 439150 -1492
rect 439218 -1548 439274 -1492
rect 439342 -1548 439398 -1492
rect 453250 4294 453306 4350
rect 453374 4294 453430 4350
rect 453498 4294 453554 4350
rect 453622 4294 453678 4350
rect 453250 4170 453306 4226
rect 453374 4170 453430 4226
rect 453498 4170 453554 4226
rect 453622 4170 453678 4226
rect 453250 4046 453306 4102
rect 453374 4046 453430 4102
rect 453498 4046 453554 4102
rect 453622 4046 453678 4102
rect 453250 3922 453306 3978
rect 453374 3922 453430 3978
rect 453498 3922 453554 3978
rect 453622 3922 453678 3978
rect 453250 -216 453306 -160
rect 453374 -216 453430 -160
rect 453498 -216 453554 -160
rect 453622 -216 453678 -160
rect 453250 -340 453306 -284
rect 453374 -340 453430 -284
rect 453498 -340 453554 -284
rect 453622 -340 453678 -284
rect 453250 -464 453306 -408
rect 453374 -464 453430 -408
rect 453498 -464 453554 -408
rect 453622 -464 453678 -408
rect 453250 -588 453306 -532
rect 453374 -588 453430 -532
rect 453498 -588 453554 -532
rect 453622 -588 453678 -532
rect 456970 10294 457026 10350
rect 457094 10294 457150 10350
rect 457218 10294 457274 10350
rect 457342 10294 457398 10350
rect 456970 10170 457026 10226
rect 457094 10170 457150 10226
rect 457218 10170 457274 10226
rect 457342 10170 457398 10226
rect 456970 10046 457026 10102
rect 457094 10046 457150 10102
rect 457218 10046 457274 10102
rect 457342 10046 457398 10102
rect 456970 9922 457026 9978
rect 457094 9922 457150 9978
rect 457218 9922 457274 9978
rect 457342 9922 457398 9978
rect 456970 -1176 457026 -1120
rect 457094 -1176 457150 -1120
rect 457218 -1176 457274 -1120
rect 457342 -1176 457398 -1120
rect 456970 -1300 457026 -1244
rect 457094 -1300 457150 -1244
rect 457218 -1300 457274 -1244
rect 457342 -1300 457398 -1244
rect 456970 -1424 457026 -1368
rect 457094 -1424 457150 -1368
rect 457218 -1424 457274 -1368
rect 457342 -1424 457398 -1368
rect 456970 -1548 457026 -1492
rect 457094 -1548 457150 -1492
rect 457218 -1548 457274 -1492
rect 457342 -1548 457398 -1492
rect 471250 4294 471306 4350
rect 471374 4294 471430 4350
rect 471498 4294 471554 4350
rect 471622 4294 471678 4350
rect 471250 4170 471306 4226
rect 471374 4170 471430 4226
rect 471498 4170 471554 4226
rect 471622 4170 471678 4226
rect 471250 4046 471306 4102
rect 471374 4046 471430 4102
rect 471498 4046 471554 4102
rect 471622 4046 471678 4102
rect 471250 3922 471306 3978
rect 471374 3922 471430 3978
rect 471498 3922 471554 3978
rect 471622 3922 471678 3978
rect 471250 -216 471306 -160
rect 471374 -216 471430 -160
rect 471498 -216 471554 -160
rect 471622 -216 471678 -160
rect 471250 -340 471306 -284
rect 471374 -340 471430 -284
rect 471498 -340 471554 -284
rect 471622 -340 471678 -284
rect 471250 -464 471306 -408
rect 471374 -464 471430 -408
rect 471498 -464 471554 -408
rect 471622 -464 471678 -408
rect 471250 -588 471306 -532
rect 471374 -588 471430 -532
rect 471498 -588 471554 -532
rect 471622 -588 471678 -532
rect 474970 10294 475026 10350
rect 475094 10294 475150 10350
rect 475218 10294 475274 10350
rect 475342 10294 475398 10350
rect 474970 10170 475026 10226
rect 475094 10170 475150 10226
rect 475218 10170 475274 10226
rect 475342 10170 475398 10226
rect 474970 10046 475026 10102
rect 475094 10046 475150 10102
rect 475218 10046 475274 10102
rect 475342 10046 475398 10102
rect 474970 9922 475026 9978
rect 475094 9922 475150 9978
rect 475218 9922 475274 9978
rect 475342 9922 475398 9978
rect 474970 -1176 475026 -1120
rect 475094 -1176 475150 -1120
rect 475218 -1176 475274 -1120
rect 475342 -1176 475398 -1120
rect 474970 -1300 475026 -1244
rect 475094 -1300 475150 -1244
rect 475218 -1300 475274 -1244
rect 475342 -1300 475398 -1244
rect 474970 -1424 475026 -1368
rect 475094 -1424 475150 -1368
rect 475218 -1424 475274 -1368
rect 475342 -1424 475398 -1368
rect 474970 -1548 475026 -1492
rect 475094 -1548 475150 -1492
rect 475218 -1548 475274 -1492
rect 475342 -1548 475398 -1492
rect 489250 4294 489306 4350
rect 489374 4294 489430 4350
rect 489498 4294 489554 4350
rect 489622 4294 489678 4350
rect 489250 4170 489306 4226
rect 489374 4170 489430 4226
rect 489498 4170 489554 4226
rect 489622 4170 489678 4226
rect 489250 4046 489306 4102
rect 489374 4046 489430 4102
rect 489498 4046 489554 4102
rect 489622 4046 489678 4102
rect 489250 3922 489306 3978
rect 489374 3922 489430 3978
rect 489498 3922 489554 3978
rect 489622 3922 489678 3978
rect 489250 -216 489306 -160
rect 489374 -216 489430 -160
rect 489498 -216 489554 -160
rect 489622 -216 489678 -160
rect 489250 -340 489306 -284
rect 489374 -340 489430 -284
rect 489498 -340 489554 -284
rect 489622 -340 489678 -284
rect 489250 -464 489306 -408
rect 489374 -464 489430 -408
rect 489498 -464 489554 -408
rect 489622 -464 489678 -408
rect 489250 -588 489306 -532
rect 489374 -588 489430 -532
rect 489498 -588 489554 -532
rect 489622 -588 489678 -532
rect 492970 10294 493026 10350
rect 493094 10294 493150 10350
rect 493218 10294 493274 10350
rect 493342 10294 493398 10350
rect 492970 10170 493026 10226
rect 493094 10170 493150 10226
rect 493218 10170 493274 10226
rect 493342 10170 493398 10226
rect 492970 10046 493026 10102
rect 493094 10046 493150 10102
rect 493218 10046 493274 10102
rect 493342 10046 493398 10102
rect 492970 9922 493026 9978
rect 493094 9922 493150 9978
rect 493218 9922 493274 9978
rect 493342 9922 493398 9978
rect 492970 -1176 493026 -1120
rect 493094 -1176 493150 -1120
rect 493218 -1176 493274 -1120
rect 493342 -1176 493398 -1120
rect 492970 -1300 493026 -1244
rect 493094 -1300 493150 -1244
rect 493218 -1300 493274 -1244
rect 493342 -1300 493398 -1244
rect 492970 -1424 493026 -1368
rect 493094 -1424 493150 -1368
rect 493218 -1424 493274 -1368
rect 493342 -1424 493398 -1368
rect 492970 -1548 493026 -1492
rect 493094 -1548 493150 -1492
rect 493218 -1548 493274 -1492
rect 493342 -1548 493398 -1492
rect 507250 4294 507306 4350
rect 507374 4294 507430 4350
rect 507498 4294 507554 4350
rect 507622 4294 507678 4350
rect 507250 4170 507306 4226
rect 507374 4170 507430 4226
rect 507498 4170 507554 4226
rect 507622 4170 507678 4226
rect 507250 4046 507306 4102
rect 507374 4046 507430 4102
rect 507498 4046 507554 4102
rect 507622 4046 507678 4102
rect 507250 3922 507306 3978
rect 507374 3922 507430 3978
rect 507498 3922 507554 3978
rect 507622 3922 507678 3978
rect 507250 -216 507306 -160
rect 507374 -216 507430 -160
rect 507498 -216 507554 -160
rect 507622 -216 507678 -160
rect 507250 -340 507306 -284
rect 507374 -340 507430 -284
rect 507498 -340 507554 -284
rect 507622 -340 507678 -284
rect 507250 -464 507306 -408
rect 507374 -464 507430 -408
rect 507498 -464 507554 -408
rect 507622 -464 507678 -408
rect 507250 -588 507306 -532
rect 507374 -588 507430 -532
rect 507498 -588 507554 -532
rect 507622 -588 507678 -532
rect 510970 10294 511026 10350
rect 511094 10294 511150 10350
rect 511218 10294 511274 10350
rect 511342 10294 511398 10350
rect 510970 10170 511026 10226
rect 511094 10170 511150 10226
rect 511218 10170 511274 10226
rect 511342 10170 511398 10226
rect 510970 10046 511026 10102
rect 511094 10046 511150 10102
rect 511218 10046 511274 10102
rect 511342 10046 511398 10102
rect 510970 9922 511026 9978
rect 511094 9922 511150 9978
rect 511218 9922 511274 9978
rect 511342 9922 511398 9978
rect 510970 -1176 511026 -1120
rect 511094 -1176 511150 -1120
rect 511218 -1176 511274 -1120
rect 511342 -1176 511398 -1120
rect 510970 -1300 511026 -1244
rect 511094 -1300 511150 -1244
rect 511218 -1300 511274 -1244
rect 511342 -1300 511398 -1244
rect 510970 -1424 511026 -1368
rect 511094 -1424 511150 -1368
rect 511218 -1424 511274 -1368
rect 511342 -1424 511398 -1368
rect 510970 -1548 511026 -1492
rect 511094 -1548 511150 -1492
rect 511218 -1548 511274 -1492
rect 511342 -1548 511398 -1492
rect 525250 4294 525306 4350
rect 525374 4294 525430 4350
rect 525498 4294 525554 4350
rect 525622 4294 525678 4350
rect 525250 4170 525306 4226
rect 525374 4170 525430 4226
rect 525498 4170 525554 4226
rect 525622 4170 525678 4226
rect 525250 4046 525306 4102
rect 525374 4046 525430 4102
rect 525498 4046 525554 4102
rect 525622 4046 525678 4102
rect 525250 3922 525306 3978
rect 525374 3922 525430 3978
rect 525498 3922 525554 3978
rect 525622 3922 525678 3978
rect 525250 -216 525306 -160
rect 525374 -216 525430 -160
rect 525498 -216 525554 -160
rect 525622 -216 525678 -160
rect 525250 -340 525306 -284
rect 525374 -340 525430 -284
rect 525498 -340 525554 -284
rect 525622 -340 525678 -284
rect 525250 -464 525306 -408
rect 525374 -464 525430 -408
rect 525498 -464 525554 -408
rect 525622 -464 525678 -408
rect 525250 -588 525306 -532
rect 525374 -588 525430 -532
rect 525498 -588 525554 -532
rect 525622 -588 525678 -532
rect 528970 598116 529026 598172
rect 529094 598116 529150 598172
rect 529218 598116 529274 598172
rect 529342 598116 529398 598172
rect 528970 597992 529026 598048
rect 529094 597992 529150 598048
rect 529218 597992 529274 598048
rect 529342 597992 529398 598048
rect 528970 597868 529026 597924
rect 529094 597868 529150 597924
rect 529218 597868 529274 597924
rect 529342 597868 529398 597924
rect 528970 597744 529026 597800
rect 529094 597744 529150 597800
rect 529218 597744 529274 597800
rect 529342 597744 529398 597800
rect 528970 586294 529026 586350
rect 529094 586294 529150 586350
rect 529218 586294 529274 586350
rect 529342 586294 529398 586350
rect 528970 586170 529026 586226
rect 529094 586170 529150 586226
rect 529218 586170 529274 586226
rect 529342 586170 529398 586226
rect 528970 586046 529026 586102
rect 529094 586046 529150 586102
rect 529218 586046 529274 586102
rect 529342 586046 529398 586102
rect 528970 585922 529026 585978
rect 529094 585922 529150 585978
rect 529218 585922 529274 585978
rect 529342 585922 529398 585978
rect 528970 568294 529026 568350
rect 529094 568294 529150 568350
rect 529218 568294 529274 568350
rect 529342 568294 529398 568350
rect 528970 568170 529026 568226
rect 529094 568170 529150 568226
rect 529218 568170 529274 568226
rect 529342 568170 529398 568226
rect 528970 568046 529026 568102
rect 529094 568046 529150 568102
rect 529218 568046 529274 568102
rect 529342 568046 529398 568102
rect 528970 567922 529026 567978
rect 529094 567922 529150 567978
rect 529218 567922 529274 567978
rect 529342 567922 529398 567978
rect 528970 550294 529026 550350
rect 529094 550294 529150 550350
rect 529218 550294 529274 550350
rect 529342 550294 529398 550350
rect 528970 550170 529026 550226
rect 529094 550170 529150 550226
rect 529218 550170 529274 550226
rect 529342 550170 529398 550226
rect 528970 550046 529026 550102
rect 529094 550046 529150 550102
rect 529218 550046 529274 550102
rect 529342 550046 529398 550102
rect 528970 549922 529026 549978
rect 529094 549922 529150 549978
rect 529218 549922 529274 549978
rect 529342 549922 529398 549978
rect 528970 532294 529026 532350
rect 529094 532294 529150 532350
rect 529218 532294 529274 532350
rect 529342 532294 529398 532350
rect 528970 532170 529026 532226
rect 529094 532170 529150 532226
rect 529218 532170 529274 532226
rect 529342 532170 529398 532226
rect 528970 532046 529026 532102
rect 529094 532046 529150 532102
rect 529218 532046 529274 532102
rect 529342 532046 529398 532102
rect 528970 531922 529026 531978
rect 529094 531922 529150 531978
rect 529218 531922 529274 531978
rect 529342 531922 529398 531978
rect 528970 514294 529026 514350
rect 529094 514294 529150 514350
rect 529218 514294 529274 514350
rect 529342 514294 529398 514350
rect 528970 514170 529026 514226
rect 529094 514170 529150 514226
rect 529218 514170 529274 514226
rect 529342 514170 529398 514226
rect 528970 514046 529026 514102
rect 529094 514046 529150 514102
rect 529218 514046 529274 514102
rect 529342 514046 529398 514102
rect 528970 513922 529026 513978
rect 529094 513922 529150 513978
rect 529218 513922 529274 513978
rect 529342 513922 529398 513978
rect 528970 496294 529026 496350
rect 529094 496294 529150 496350
rect 529218 496294 529274 496350
rect 529342 496294 529398 496350
rect 528970 496170 529026 496226
rect 529094 496170 529150 496226
rect 529218 496170 529274 496226
rect 529342 496170 529398 496226
rect 528970 496046 529026 496102
rect 529094 496046 529150 496102
rect 529218 496046 529274 496102
rect 529342 496046 529398 496102
rect 528970 495922 529026 495978
rect 529094 495922 529150 495978
rect 529218 495922 529274 495978
rect 529342 495922 529398 495978
rect 528970 478294 529026 478350
rect 529094 478294 529150 478350
rect 529218 478294 529274 478350
rect 529342 478294 529398 478350
rect 528970 478170 529026 478226
rect 529094 478170 529150 478226
rect 529218 478170 529274 478226
rect 529342 478170 529398 478226
rect 528970 478046 529026 478102
rect 529094 478046 529150 478102
rect 529218 478046 529274 478102
rect 529342 478046 529398 478102
rect 528970 477922 529026 477978
rect 529094 477922 529150 477978
rect 529218 477922 529274 477978
rect 529342 477922 529398 477978
rect 528970 460294 529026 460350
rect 529094 460294 529150 460350
rect 529218 460294 529274 460350
rect 529342 460294 529398 460350
rect 528970 460170 529026 460226
rect 529094 460170 529150 460226
rect 529218 460170 529274 460226
rect 529342 460170 529398 460226
rect 528970 460046 529026 460102
rect 529094 460046 529150 460102
rect 529218 460046 529274 460102
rect 529342 460046 529398 460102
rect 528970 459922 529026 459978
rect 529094 459922 529150 459978
rect 529218 459922 529274 459978
rect 529342 459922 529398 459978
rect 528970 442294 529026 442350
rect 529094 442294 529150 442350
rect 529218 442294 529274 442350
rect 529342 442294 529398 442350
rect 528970 442170 529026 442226
rect 529094 442170 529150 442226
rect 529218 442170 529274 442226
rect 529342 442170 529398 442226
rect 528970 442046 529026 442102
rect 529094 442046 529150 442102
rect 529218 442046 529274 442102
rect 529342 442046 529398 442102
rect 528970 441922 529026 441978
rect 529094 441922 529150 441978
rect 529218 441922 529274 441978
rect 529342 441922 529398 441978
rect 528970 424294 529026 424350
rect 529094 424294 529150 424350
rect 529218 424294 529274 424350
rect 529342 424294 529398 424350
rect 528970 424170 529026 424226
rect 529094 424170 529150 424226
rect 529218 424170 529274 424226
rect 529342 424170 529398 424226
rect 528970 424046 529026 424102
rect 529094 424046 529150 424102
rect 529218 424046 529274 424102
rect 529342 424046 529398 424102
rect 528970 423922 529026 423978
rect 529094 423922 529150 423978
rect 529218 423922 529274 423978
rect 529342 423922 529398 423978
rect 528970 406294 529026 406350
rect 529094 406294 529150 406350
rect 529218 406294 529274 406350
rect 529342 406294 529398 406350
rect 528970 406170 529026 406226
rect 529094 406170 529150 406226
rect 529218 406170 529274 406226
rect 529342 406170 529398 406226
rect 528970 406046 529026 406102
rect 529094 406046 529150 406102
rect 529218 406046 529274 406102
rect 529342 406046 529398 406102
rect 528970 405922 529026 405978
rect 529094 405922 529150 405978
rect 529218 405922 529274 405978
rect 529342 405922 529398 405978
rect 528970 388294 529026 388350
rect 529094 388294 529150 388350
rect 529218 388294 529274 388350
rect 529342 388294 529398 388350
rect 528970 388170 529026 388226
rect 529094 388170 529150 388226
rect 529218 388170 529274 388226
rect 529342 388170 529398 388226
rect 528970 388046 529026 388102
rect 529094 388046 529150 388102
rect 529218 388046 529274 388102
rect 529342 388046 529398 388102
rect 528970 387922 529026 387978
rect 529094 387922 529150 387978
rect 529218 387922 529274 387978
rect 529342 387922 529398 387978
rect 528970 370294 529026 370350
rect 529094 370294 529150 370350
rect 529218 370294 529274 370350
rect 529342 370294 529398 370350
rect 528970 370170 529026 370226
rect 529094 370170 529150 370226
rect 529218 370170 529274 370226
rect 529342 370170 529398 370226
rect 528970 370046 529026 370102
rect 529094 370046 529150 370102
rect 529218 370046 529274 370102
rect 529342 370046 529398 370102
rect 528970 369922 529026 369978
rect 529094 369922 529150 369978
rect 529218 369922 529274 369978
rect 529342 369922 529398 369978
rect 528970 352294 529026 352350
rect 529094 352294 529150 352350
rect 529218 352294 529274 352350
rect 529342 352294 529398 352350
rect 528970 352170 529026 352226
rect 529094 352170 529150 352226
rect 529218 352170 529274 352226
rect 529342 352170 529398 352226
rect 528970 352046 529026 352102
rect 529094 352046 529150 352102
rect 529218 352046 529274 352102
rect 529342 352046 529398 352102
rect 528970 351922 529026 351978
rect 529094 351922 529150 351978
rect 529218 351922 529274 351978
rect 529342 351922 529398 351978
rect 528970 334294 529026 334350
rect 529094 334294 529150 334350
rect 529218 334294 529274 334350
rect 529342 334294 529398 334350
rect 528970 334170 529026 334226
rect 529094 334170 529150 334226
rect 529218 334170 529274 334226
rect 529342 334170 529398 334226
rect 528970 334046 529026 334102
rect 529094 334046 529150 334102
rect 529218 334046 529274 334102
rect 529342 334046 529398 334102
rect 528970 333922 529026 333978
rect 529094 333922 529150 333978
rect 529218 333922 529274 333978
rect 529342 333922 529398 333978
rect 528970 316294 529026 316350
rect 529094 316294 529150 316350
rect 529218 316294 529274 316350
rect 529342 316294 529398 316350
rect 528970 316170 529026 316226
rect 529094 316170 529150 316226
rect 529218 316170 529274 316226
rect 529342 316170 529398 316226
rect 528970 316046 529026 316102
rect 529094 316046 529150 316102
rect 529218 316046 529274 316102
rect 529342 316046 529398 316102
rect 528970 315922 529026 315978
rect 529094 315922 529150 315978
rect 529218 315922 529274 315978
rect 529342 315922 529398 315978
rect 528970 298294 529026 298350
rect 529094 298294 529150 298350
rect 529218 298294 529274 298350
rect 529342 298294 529398 298350
rect 528970 298170 529026 298226
rect 529094 298170 529150 298226
rect 529218 298170 529274 298226
rect 529342 298170 529398 298226
rect 528970 298046 529026 298102
rect 529094 298046 529150 298102
rect 529218 298046 529274 298102
rect 529342 298046 529398 298102
rect 528970 297922 529026 297978
rect 529094 297922 529150 297978
rect 529218 297922 529274 297978
rect 529342 297922 529398 297978
rect 528970 280294 529026 280350
rect 529094 280294 529150 280350
rect 529218 280294 529274 280350
rect 529342 280294 529398 280350
rect 528970 280170 529026 280226
rect 529094 280170 529150 280226
rect 529218 280170 529274 280226
rect 529342 280170 529398 280226
rect 528970 280046 529026 280102
rect 529094 280046 529150 280102
rect 529218 280046 529274 280102
rect 529342 280046 529398 280102
rect 528970 279922 529026 279978
rect 529094 279922 529150 279978
rect 529218 279922 529274 279978
rect 529342 279922 529398 279978
rect 528970 262294 529026 262350
rect 529094 262294 529150 262350
rect 529218 262294 529274 262350
rect 529342 262294 529398 262350
rect 528970 262170 529026 262226
rect 529094 262170 529150 262226
rect 529218 262170 529274 262226
rect 529342 262170 529398 262226
rect 528970 262046 529026 262102
rect 529094 262046 529150 262102
rect 529218 262046 529274 262102
rect 529342 262046 529398 262102
rect 528970 261922 529026 261978
rect 529094 261922 529150 261978
rect 529218 261922 529274 261978
rect 529342 261922 529398 261978
rect 528970 244294 529026 244350
rect 529094 244294 529150 244350
rect 529218 244294 529274 244350
rect 529342 244294 529398 244350
rect 528970 244170 529026 244226
rect 529094 244170 529150 244226
rect 529218 244170 529274 244226
rect 529342 244170 529398 244226
rect 528970 244046 529026 244102
rect 529094 244046 529150 244102
rect 529218 244046 529274 244102
rect 529342 244046 529398 244102
rect 528970 243922 529026 243978
rect 529094 243922 529150 243978
rect 529218 243922 529274 243978
rect 529342 243922 529398 243978
rect 528970 226294 529026 226350
rect 529094 226294 529150 226350
rect 529218 226294 529274 226350
rect 529342 226294 529398 226350
rect 528970 226170 529026 226226
rect 529094 226170 529150 226226
rect 529218 226170 529274 226226
rect 529342 226170 529398 226226
rect 528970 226046 529026 226102
rect 529094 226046 529150 226102
rect 529218 226046 529274 226102
rect 529342 226046 529398 226102
rect 528970 225922 529026 225978
rect 529094 225922 529150 225978
rect 529218 225922 529274 225978
rect 529342 225922 529398 225978
rect 528970 208294 529026 208350
rect 529094 208294 529150 208350
rect 529218 208294 529274 208350
rect 529342 208294 529398 208350
rect 528970 208170 529026 208226
rect 529094 208170 529150 208226
rect 529218 208170 529274 208226
rect 529342 208170 529398 208226
rect 528970 208046 529026 208102
rect 529094 208046 529150 208102
rect 529218 208046 529274 208102
rect 529342 208046 529398 208102
rect 528970 207922 529026 207978
rect 529094 207922 529150 207978
rect 529218 207922 529274 207978
rect 529342 207922 529398 207978
rect 528970 190294 529026 190350
rect 529094 190294 529150 190350
rect 529218 190294 529274 190350
rect 529342 190294 529398 190350
rect 528970 190170 529026 190226
rect 529094 190170 529150 190226
rect 529218 190170 529274 190226
rect 529342 190170 529398 190226
rect 528970 190046 529026 190102
rect 529094 190046 529150 190102
rect 529218 190046 529274 190102
rect 529342 190046 529398 190102
rect 528970 189922 529026 189978
rect 529094 189922 529150 189978
rect 529218 189922 529274 189978
rect 529342 189922 529398 189978
rect 528970 172294 529026 172350
rect 529094 172294 529150 172350
rect 529218 172294 529274 172350
rect 529342 172294 529398 172350
rect 528970 172170 529026 172226
rect 529094 172170 529150 172226
rect 529218 172170 529274 172226
rect 529342 172170 529398 172226
rect 528970 172046 529026 172102
rect 529094 172046 529150 172102
rect 529218 172046 529274 172102
rect 529342 172046 529398 172102
rect 528970 171922 529026 171978
rect 529094 171922 529150 171978
rect 529218 171922 529274 171978
rect 529342 171922 529398 171978
rect 528970 154294 529026 154350
rect 529094 154294 529150 154350
rect 529218 154294 529274 154350
rect 529342 154294 529398 154350
rect 528970 154170 529026 154226
rect 529094 154170 529150 154226
rect 529218 154170 529274 154226
rect 529342 154170 529398 154226
rect 528970 154046 529026 154102
rect 529094 154046 529150 154102
rect 529218 154046 529274 154102
rect 529342 154046 529398 154102
rect 528970 153922 529026 153978
rect 529094 153922 529150 153978
rect 529218 153922 529274 153978
rect 529342 153922 529398 153978
rect 528970 136294 529026 136350
rect 529094 136294 529150 136350
rect 529218 136294 529274 136350
rect 529342 136294 529398 136350
rect 528970 136170 529026 136226
rect 529094 136170 529150 136226
rect 529218 136170 529274 136226
rect 529342 136170 529398 136226
rect 528970 136046 529026 136102
rect 529094 136046 529150 136102
rect 529218 136046 529274 136102
rect 529342 136046 529398 136102
rect 528970 135922 529026 135978
rect 529094 135922 529150 135978
rect 529218 135922 529274 135978
rect 529342 135922 529398 135978
rect 528970 118294 529026 118350
rect 529094 118294 529150 118350
rect 529218 118294 529274 118350
rect 529342 118294 529398 118350
rect 528970 118170 529026 118226
rect 529094 118170 529150 118226
rect 529218 118170 529274 118226
rect 529342 118170 529398 118226
rect 528970 118046 529026 118102
rect 529094 118046 529150 118102
rect 529218 118046 529274 118102
rect 529342 118046 529398 118102
rect 528970 117922 529026 117978
rect 529094 117922 529150 117978
rect 529218 117922 529274 117978
rect 529342 117922 529398 117978
rect 528970 100294 529026 100350
rect 529094 100294 529150 100350
rect 529218 100294 529274 100350
rect 529342 100294 529398 100350
rect 528970 100170 529026 100226
rect 529094 100170 529150 100226
rect 529218 100170 529274 100226
rect 529342 100170 529398 100226
rect 528970 100046 529026 100102
rect 529094 100046 529150 100102
rect 529218 100046 529274 100102
rect 529342 100046 529398 100102
rect 528970 99922 529026 99978
rect 529094 99922 529150 99978
rect 529218 99922 529274 99978
rect 529342 99922 529398 99978
rect 528970 82294 529026 82350
rect 529094 82294 529150 82350
rect 529218 82294 529274 82350
rect 529342 82294 529398 82350
rect 528970 82170 529026 82226
rect 529094 82170 529150 82226
rect 529218 82170 529274 82226
rect 529342 82170 529398 82226
rect 528970 82046 529026 82102
rect 529094 82046 529150 82102
rect 529218 82046 529274 82102
rect 529342 82046 529398 82102
rect 528970 81922 529026 81978
rect 529094 81922 529150 81978
rect 529218 81922 529274 81978
rect 529342 81922 529398 81978
rect 528970 64294 529026 64350
rect 529094 64294 529150 64350
rect 529218 64294 529274 64350
rect 529342 64294 529398 64350
rect 528970 64170 529026 64226
rect 529094 64170 529150 64226
rect 529218 64170 529274 64226
rect 529342 64170 529398 64226
rect 528970 64046 529026 64102
rect 529094 64046 529150 64102
rect 529218 64046 529274 64102
rect 529342 64046 529398 64102
rect 528970 63922 529026 63978
rect 529094 63922 529150 63978
rect 529218 63922 529274 63978
rect 529342 63922 529398 63978
rect 528970 46294 529026 46350
rect 529094 46294 529150 46350
rect 529218 46294 529274 46350
rect 529342 46294 529398 46350
rect 528970 46170 529026 46226
rect 529094 46170 529150 46226
rect 529218 46170 529274 46226
rect 529342 46170 529398 46226
rect 528970 46046 529026 46102
rect 529094 46046 529150 46102
rect 529218 46046 529274 46102
rect 529342 46046 529398 46102
rect 528970 45922 529026 45978
rect 529094 45922 529150 45978
rect 529218 45922 529274 45978
rect 529342 45922 529398 45978
rect 528970 28294 529026 28350
rect 529094 28294 529150 28350
rect 529218 28294 529274 28350
rect 529342 28294 529398 28350
rect 528970 28170 529026 28226
rect 529094 28170 529150 28226
rect 529218 28170 529274 28226
rect 529342 28170 529398 28226
rect 528970 28046 529026 28102
rect 529094 28046 529150 28102
rect 529218 28046 529274 28102
rect 529342 28046 529398 28102
rect 528970 27922 529026 27978
rect 529094 27922 529150 27978
rect 529218 27922 529274 27978
rect 529342 27922 529398 27978
rect 528970 10294 529026 10350
rect 529094 10294 529150 10350
rect 529218 10294 529274 10350
rect 529342 10294 529398 10350
rect 528970 10170 529026 10226
rect 529094 10170 529150 10226
rect 529218 10170 529274 10226
rect 529342 10170 529398 10226
rect 528970 10046 529026 10102
rect 529094 10046 529150 10102
rect 529218 10046 529274 10102
rect 529342 10046 529398 10102
rect 528970 9922 529026 9978
rect 529094 9922 529150 9978
rect 529218 9922 529274 9978
rect 529342 9922 529398 9978
rect 528970 -1176 529026 -1120
rect 529094 -1176 529150 -1120
rect 529218 -1176 529274 -1120
rect 529342 -1176 529398 -1120
rect 528970 -1300 529026 -1244
rect 529094 -1300 529150 -1244
rect 529218 -1300 529274 -1244
rect 529342 -1300 529398 -1244
rect 528970 -1424 529026 -1368
rect 529094 -1424 529150 -1368
rect 529218 -1424 529274 -1368
rect 529342 -1424 529398 -1368
rect 528970 -1548 529026 -1492
rect 529094 -1548 529150 -1492
rect 529218 -1548 529274 -1492
rect 529342 -1548 529398 -1492
rect 543250 597156 543306 597212
rect 543374 597156 543430 597212
rect 543498 597156 543554 597212
rect 543622 597156 543678 597212
rect 543250 597032 543306 597088
rect 543374 597032 543430 597088
rect 543498 597032 543554 597088
rect 543622 597032 543678 597088
rect 543250 596908 543306 596964
rect 543374 596908 543430 596964
rect 543498 596908 543554 596964
rect 543622 596908 543678 596964
rect 543250 596784 543306 596840
rect 543374 596784 543430 596840
rect 543498 596784 543554 596840
rect 543622 596784 543678 596840
rect 543250 580294 543306 580350
rect 543374 580294 543430 580350
rect 543498 580294 543554 580350
rect 543622 580294 543678 580350
rect 543250 580170 543306 580226
rect 543374 580170 543430 580226
rect 543498 580170 543554 580226
rect 543622 580170 543678 580226
rect 543250 580046 543306 580102
rect 543374 580046 543430 580102
rect 543498 580046 543554 580102
rect 543622 580046 543678 580102
rect 543250 579922 543306 579978
rect 543374 579922 543430 579978
rect 543498 579922 543554 579978
rect 543622 579922 543678 579978
rect 543250 562294 543306 562350
rect 543374 562294 543430 562350
rect 543498 562294 543554 562350
rect 543622 562294 543678 562350
rect 543250 562170 543306 562226
rect 543374 562170 543430 562226
rect 543498 562170 543554 562226
rect 543622 562170 543678 562226
rect 543250 562046 543306 562102
rect 543374 562046 543430 562102
rect 543498 562046 543554 562102
rect 543622 562046 543678 562102
rect 543250 561922 543306 561978
rect 543374 561922 543430 561978
rect 543498 561922 543554 561978
rect 543622 561922 543678 561978
rect 543250 544294 543306 544350
rect 543374 544294 543430 544350
rect 543498 544294 543554 544350
rect 543622 544294 543678 544350
rect 543250 544170 543306 544226
rect 543374 544170 543430 544226
rect 543498 544170 543554 544226
rect 543622 544170 543678 544226
rect 543250 544046 543306 544102
rect 543374 544046 543430 544102
rect 543498 544046 543554 544102
rect 543622 544046 543678 544102
rect 543250 543922 543306 543978
rect 543374 543922 543430 543978
rect 543498 543922 543554 543978
rect 543622 543922 543678 543978
rect 543250 526294 543306 526350
rect 543374 526294 543430 526350
rect 543498 526294 543554 526350
rect 543622 526294 543678 526350
rect 543250 526170 543306 526226
rect 543374 526170 543430 526226
rect 543498 526170 543554 526226
rect 543622 526170 543678 526226
rect 543250 526046 543306 526102
rect 543374 526046 543430 526102
rect 543498 526046 543554 526102
rect 543622 526046 543678 526102
rect 543250 525922 543306 525978
rect 543374 525922 543430 525978
rect 543498 525922 543554 525978
rect 543622 525922 543678 525978
rect 543250 508294 543306 508350
rect 543374 508294 543430 508350
rect 543498 508294 543554 508350
rect 543622 508294 543678 508350
rect 543250 508170 543306 508226
rect 543374 508170 543430 508226
rect 543498 508170 543554 508226
rect 543622 508170 543678 508226
rect 543250 508046 543306 508102
rect 543374 508046 543430 508102
rect 543498 508046 543554 508102
rect 543622 508046 543678 508102
rect 543250 507922 543306 507978
rect 543374 507922 543430 507978
rect 543498 507922 543554 507978
rect 543622 507922 543678 507978
rect 543250 490294 543306 490350
rect 543374 490294 543430 490350
rect 543498 490294 543554 490350
rect 543622 490294 543678 490350
rect 543250 490170 543306 490226
rect 543374 490170 543430 490226
rect 543498 490170 543554 490226
rect 543622 490170 543678 490226
rect 543250 490046 543306 490102
rect 543374 490046 543430 490102
rect 543498 490046 543554 490102
rect 543622 490046 543678 490102
rect 543250 489922 543306 489978
rect 543374 489922 543430 489978
rect 543498 489922 543554 489978
rect 543622 489922 543678 489978
rect 543250 472294 543306 472350
rect 543374 472294 543430 472350
rect 543498 472294 543554 472350
rect 543622 472294 543678 472350
rect 543250 472170 543306 472226
rect 543374 472170 543430 472226
rect 543498 472170 543554 472226
rect 543622 472170 543678 472226
rect 543250 472046 543306 472102
rect 543374 472046 543430 472102
rect 543498 472046 543554 472102
rect 543622 472046 543678 472102
rect 543250 471922 543306 471978
rect 543374 471922 543430 471978
rect 543498 471922 543554 471978
rect 543622 471922 543678 471978
rect 543250 454294 543306 454350
rect 543374 454294 543430 454350
rect 543498 454294 543554 454350
rect 543622 454294 543678 454350
rect 543250 454170 543306 454226
rect 543374 454170 543430 454226
rect 543498 454170 543554 454226
rect 543622 454170 543678 454226
rect 543250 454046 543306 454102
rect 543374 454046 543430 454102
rect 543498 454046 543554 454102
rect 543622 454046 543678 454102
rect 543250 453922 543306 453978
rect 543374 453922 543430 453978
rect 543498 453922 543554 453978
rect 543622 453922 543678 453978
rect 543250 436294 543306 436350
rect 543374 436294 543430 436350
rect 543498 436294 543554 436350
rect 543622 436294 543678 436350
rect 543250 436170 543306 436226
rect 543374 436170 543430 436226
rect 543498 436170 543554 436226
rect 543622 436170 543678 436226
rect 543250 436046 543306 436102
rect 543374 436046 543430 436102
rect 543498 436046 543554 436102
rect 543622 436046 543678 436102
rect 543250 435922 543306 435978
rect 543374 435922 543430 435978
rect 543498 435922 543554 435978
rect 543622 435922 543678 435978
rect 543250 418294 543306 418350
rect 543374 418294 543430 418350
rect 543498 418294 543554 418350
rect 543622 418294 543678 418350
rect 543250 418170 543306 418226
rect 543374 418170 543430 418226
rect 543498 418170 543554 418226
rect 543622 418170 543678 418226
rect 543250 418046 543306 418102
rect 543374 418046 543430 418102
rect 543498 418046 543554 418102
rect 543622 418046 543678 418102
rect 543250 417922 543306 417978
rect 543374 417922 543430 417978
rect 543498 417922 543554 417978
rect 543622 417922 543678 417978
rect 543250 400294 543306 400350
rect 543374 400294 543430 400350
rect 543498 400294 543554 400350
rect 543622 400294 543678 400350
rect 543250 400170 543306 400226
rect 543374 400170 543430 400226
rect 543498 400170 543554 400226
rect 543622 400170 543678 400226
rect 543250 400046 543306 400102
rect 543374 400046 543430 400102
rect 543498 400046 543554 400102
rect 543622 400046 543678 400102
rect 543250 399922 543306 399978
rect 543374 399922 543430 399978
rect 543498 399922 543554 399978
rect 543622 399922 543678 399978
rect 543250 382294 543306 382350
rect 543374 382294 543430 382350
rect 543498 382294 543554 382350
rect 543622 382294 543678 382350
rect 543250 382170 543306 382226
rect 543374 382170 543430 382226
rect 543498 382170 543554 382226
rect 543622 382170 543678 382226
rect 543250 382046 543306 382102
rect 543374 382046 543430 382102
rect 543498 382046 543554 382102
rect 543622 382046 543678 382102
rect 543250 381922 543306 381978
rect 543374 381922 543430 381978
rect 543498 381922 543554 381978
rect 543622 381922 543678 381978
rect 543250 364294 543306 364350
rect 543374 364294 543430 364350
rect 543498 364294 543554 364350
rect 543622 364294 543678 364350
rect 543250 364170 543306 364226
rect 543374 364170 543430 364226
rect 543498 364170 543554 364226
rect 543622 364170 543678 364226
rect 543250 364046 543306 364102
rect 543374 364046 543430 364102
rect 543498 364046 543554 364102
rect 543622 364046 543678 364102
rect 543250 363922 543306 363978
rect 543374 363922 543430 363978
rect 543498 363922 543554 363978
rect 543622 363922 543678 363978
rect 543250 346294 543306 346350
rect 543374 346294 543430 346350
rect 543498 346294 543554 346350
rect 543622 346294 543678 346350
rect 543250 346170 543306 346226
rect 543374 346170 543430 346226
rect 543498 346170 543554 346226
rect 543622 346170 543678 346226
rect 543250 346046 543306 346102
rect 543374 346046 543430 346102
rect 543498 346046 543554 346102
rect 543622 346046 543678 346102
rect 543250 345922 543306 345978
rect 543374 345922 543430 345978
rect 543498 345922 543554 345978
rect 543622 345922 543678 345978
rect 543250 328294 543306 328350
rect 543374 328294 543430 328350
rect 543498 328294 543554 328350
rect 543622 328294 543678 328350
rect 543250 328170 543306 328226
rect 543374 328170 543430 328226
rect 543498 328170 543554 328226
rect 543622 328170 543678 328226
rect 543250 328046 543306 328102
rect 543374 328046 543430 328102
rect 543498 328046 543554 328102
rect 543622 328046 543678 328102
rect 543250 327922 543306 327978
rect 543374 327922 543430 327978
rect 543498 327922 543554 327978
rect 543622 327922 543678 327978
rect 543250 310294 543306 310350
rect 543374 310294 543430 310350
rect 543498 310294 543554 310350
rect 543622 310294 543678 310350
rect 543250 310170 543306 310226
rect 543374 310170 543430 310226
rect 543498 310170 543554 310226
rect 543622 310170 543678 310226
rect 543250 310046 543306 310102
rect 543374 310046 543430 310102
rect 543498 310046 543554 310102
rect 543622 310046 543678 310102
rect 543250 309922 543306 309978
rect 543374 309922 543430 309978
rect 543498 309922 543554 309978
rect 543622 309922 543678 309978
rect 543250 292294 543306 292350
rect 543374 292294 543430 292350
rect 543498 292294 543554 292350
rect 543622 292294 543678 292350
rect 543250 292170 543306 292226
rect 543374 292170 543430 292226
rect 543498 292170 543554 292226
rect 543622 292170 543678 292226
rect 543250 292046 543306 292102
rect 543374 292046 543430 292102
rect 543498 292046 543554 292102
rect 543622 292046 543678 292102
rect 543250 291922 543306 291978
rect 543374 291922 543430 291978
rect 543498 291922 543554 291978
rect 543622 291922 543678 291978
rect 543250 274294 543306 274350
rect 543374 274294 543430 274350
rect 543498 274294 543554 274350
rect 543622 274294 543678 274350
rect 543250 274170 543306 274226
rect 543374 274170 543430 274226
rect 543498 274170 543554 274226
rect 543622 274170 543678 274226
rect 543250 274046 543306 274102
rect 543374 274046 543430 274102
rect 543498 274046 543554 274102
rect 543622 274046 543678 274102
rect 543250 273922 543306 273978
rect 543374 273922 543430 273978
rect 543498 273922 543554 273978
rect 543622 273922 543678 273978
rect 543250 256294 543306 256350
rect 543374 256294 543430 256350
rect 543498 256294 543554 256350
rect 543622 256294 543678 256350
rect 543250 256170 543306 256226
rect 543374 256170 543430 256226
rect 543498 256170 543554 256226
rect 543622 256170 543678 256226
rect 543250 256046 543306 256102
rect 543374 256046 543430 256102
rect 543498 256046 543554 256102
rect 543622 256046 543678 256102
rect 543250 255922 543306 255978
rect 543374 255922 543430 255978
rect 543498 255922 543554 255978
rect 543622 255922 543678 255978
rect 543250 238294 543306 238350
rect 543374 238294 543430 238350
rect 543498 238294 543554 238350
rect 543622 238294 543678 238350
rect 543250 238170 543306 238226
rect 543374 238170 543430 238226
rect 543498 238170 543554 238226
rect 543622 238170 543678 238226
rect 543250 238046 543306 238102
rect 543374 238046 543430 238102
rect 543498 238046 543554 238102
rect 543622 238046 543678 238102
rect 543250 237922 543306 237978
rect 543374 237922 543430 237978
rect 543498 237922 543554 237978
rect 543622 237922 543678 237978
rect 543250 220294 543306 220350
rect 543374 220294 543430 220350
rect 543498 220294 543554 220350
rect 543622 220294 543678 220350
rect 543250 220170 543306 220226
rect 543374 220170 543430 220226
rect 543498 220170 543554 220226
rect 543622 220170 543678 220226
rect 543250 220046 543306 220102
rect 543374 220046 543430 220102
rect 543498 220046 543554 220102
rect 543622 220046 543678 220102
rect 543250 219922 543306 219978
rect 543374 219922 543430 219978
rect 543498 219922 543554 219978
rect 543622 219922 543678 219978
rect 543250 202294 543306 202350
rect 543374 202294 543430 202350
rect 543498 202294 543554 202350
rect 543622 202294 543678 202350
rect 543250 202170 543306 202226
rect 543374 202170 543430 202226
rect 543498 202170 543554 202226
rect 543622 202170 543678 202226
rect 543250 202046 543306 202102
rect 543374 202046 543430 202102
rect 543498 202046 543554 202102
rect 543622 202046 543678 202102
rect 543250 201922 543306 201978
rect 543374 201922 543430 201978
rect 543498 201922 543554 201978
rect 543622 201922 543678 201978
rect 543250 184294 543306 184350
rect 543374 184294 543430 184350
rect 543498 184294 543554 184350
rect 543622 184294 543678 184350
rect 543250 184170 543306 184226
rect 543374 184170 543430 184226
rect 543498 184170 543554 184226
rect 543622 184170 543678 184226
rect 543250 184046 543306 184102
rect 543374 184046 543430 184102
rect 543498 184046 543554 184102
rect 543622 184046 543678 184102
rect 543250 183922 543306 183978
rect 543374 183922 543430 183978
rect 543498 183922 543554 183978
rect 543622 183922 543678 183978
rect 543250 166294 543306 166350
rect 543374 166294 543430 166350
rect 543498 166294 543554 166350
rect 543622 166294 543678 166350
rect 543250 166170 543306 166226
rect 543374 166170 543430 166226
rect 543498 166170 543554 166226
rect 543622 166170 543678 166226
rect 543250 166046 543306 166102
rect 543374 166046 543430 166102
rect 543498 166046 543554 166102
rect 543622 166046 543678 166102
rect 543250 165922 543306 165978
rect 543374 165922 543430 165978
rect 543498 165922 543554 165978
rect 543622 165922 543678 165978
rect 543250 148294 543306 148350
rect 543374 148294 543430 148350
rect 543498 148294 543554 148350
rect 543622 148294 543678 148350
rect 543250 148170 543306 148226
rect 543374 148170 543430 148226
rect 543498 148170 543554 148226
rect 543622 148170 543678 148226
rect 543250 148046 543306 148102
rect 543374 148046 543430 148102
rect 543498 148046 543554 148102
rect 543622 148046 543678 148102
rect 543250 147922 543306 147978
rect 543374 147922 543430 147978
rect 543498 147922 543554 147978
rect 543622 147922 543678 147978
rect 543250 130294 543306 130350
rect 543374 130294 543430 130350
rect 543498 130294 543554 130350
rect 543622 130294 543678 130350
rect 543250 130170 543306 130226
rect 543374 130170 543430 130226
rect 543498 130170 543554 130226
rect 543622 130170 543678 130226
rect 543250 130046 543306 130102
rect 543374 130046 543430 130102
rect 543498 130046 543554 130102
rect 543622 130046 543678 130102
rect 543250 129922 543306 129978
rect 543374 129922 543430 129978
rect 543498 129922 543554 129978
rect 543622 129922 543678 129978
rect 543250 112294 543306 112350
rect 543374 112294 543430 112350
rect 543498 112294 543554 112350
rect 543622 112294 543678 112350
rect 543250 112170 543306 112226
rect 543374 112170 543430 112226
rect 543498 112170 543554 112226
rect 543622 112170 543678 112226
rect 543250 112046 543306 112102
rect 543374 112046 543430 112102
rect 543498 112046 543554 112102
rect 543622 112046 543678 112102
rect 543250 111922 543306 111978
rect 543374 111922 543430 111978
rect 543498 111922 543554 111978
rect 543622 111922 543678 111978
rect 543250 94294 543306 94350
rect 543374 94294 543430 94350
rect 543498 94294 543554 94350
rect 543622 94294 543678 94350
rect 543250 94170 543306 94226
rect 543374 94170 543430 94226
rect 543498 94170 543554 94226
rect 543622 94170 543678 94226
rect 543250 94046 543306 94102
rect 543374 94046 543430 94102
rect 543498 94046 543554 94102
rect 543622 94046 543678 94102
rect 543250 93922 543306 93978
rect 543374 93922 543430 93978
rect 543498 93922 543554 93978
rect 543622 93922 543678 93978
rect 543250 76294 543306 76350
rect 543374 76294 543430 76350
rect 543498 76294 543554 76350
rect 543622 76294 543678 76350
rect 543250 76170 543306 76226
rect 543374 76170 543430 76226
rect 543498 76170 543554 76226
rect 543622 76170 543678 76226
rect 543250 76046 543306 76102
rect 543374 76046 543430 76102
rect 543498 76046 543554 76102
rect 543622 76046 543678 76102
rect 543250 75922 543306 75978
rect 543374 75922 543430 75978
rect 543498 75922 543554 75978
rect 543622 75922 543678 75978
rect 543250 58294 543306 58350
rect 543374 58294 543430 58350
rect 543498 58294 543554 58350
rect 543622 58294 543678 58350
rect 543250 58170 543306 58226
rect 543374 58170 543430 58226
rect 543498 58170 543554 58226
rect 543622 58170 543678 58226
rect 543250 58046 543306 58102
rect 543374 58046 543430 58102
rect 543498 58046 543554 58102
rect 543622 58046 543678 58102
rect 543250 57922 543306 57978
rect 543374 57922 543430 57978
rect 543498 57922 543554 57978
rect 543622 57922 543678 57978
rect 543250 40294 543306 40350
rect 543374 40294 543430 40350
rect 543498 40294 543554 40350
rect 543622 40294 543678 40350
rect 543250 40170 543306 40226
rect 543374 40170 543430 40226
rect 543498 40170 543554 40226
rect 543622 40170 543678 40226
rect 543250 40046 543306 40102
rect 543374 40046 543430 40102
rect 543498 40046 543554 40102
rect 543622 40046 543678 40102
rect 543250 39922 543306 39978
rect 543374 39922 543430 39978
rect 543498 39922 543554 39978
rect 543622 39922 543678 39978
rect 543250 22294 543306 22350
rect 543374 22294 543430 22350
rect 543498 22294 543554 22350
rect 543622 22294 543678 22350
rect 543250 22170 543306 22226
rect 543374 22170 543430 22226
rect 543498 22170 543554 22226
rect 543622 22170 543678 22226
rect 543250 22046 543306 22102
rect 543374 22046 543430 22102
rect 543498 22046 543554 22102
rect 543622 22046 543678 22102
rect 543250 21922 543306 21978
rect 543374 21922 543430 21978
rect 543498 21922 543554 21978
rect 543622 21922 543678 21978
rect 543250 4294 543306 4350
rect 543374 4294 543430 4350
rect 543498 4294 543554 4350
rect 543622 4294 543678 4350
rect 543250 4170 543306 4226
rect 543374 4170 543430 4226
rect 543498 4170 543554 4226
rect 543622 4170 543678 4226
rect 543250 4046 543306 4102
rect 543374 4046 543430 4102
rect 543498 4046 543554 4102
rect 543622 4046 543678 4102
rect 543250 3922 543306 3978
rect 543374 3922 543430 3978
rect 543498 3922 543554 3978
rect 543622 3922 543678 3978
rect 543250 -216 543306 -160
rect 543374 -216 543430 -160
rect 543498 -216 543554 -160
rect 543622 -216 543678 -160
rect 543250 -340 543306 -284
rect 543374 -340 543430 -284
rect 543498 -340 543554 -284
rect 543622 -340 543678 -284
rect 543250 -464 543306 -408
rect 543374 -464 543430 -408
rect 543498 -464 543554 -408
rect 543622 -464 543678 -408
rect 543250 -588 543306 -532
rect 543374 -588 543430 -532
rect 543498 -588 543554 -532
rect 543622 -588 543678 -532
rect 546970 598116 547026 598172
rect 547094 598116 547150 598172
rect 547218 598116 547274 598172
rect 547342 598116 547398 598172
rect 546970 597992 547026 598048
rect 547094 597992 547150 598048
rect 547218 597992 547274 598048
rect 547342 597992 547398 598048
rect 546970 597868 547026 597924
rect 547094 597868 547150 597924
rect 547218 597868 547274 597924
rect 547342 597868 547398 597924
rect 546970 597744 547026 597800
rect 547094 597744 547150 597800
rect 547218 597744 547274 597800
rect 547342 597744 547398 597800
rect 546970 586294 547026 586350
rect 547094 586294 547150 586350
rect 547218 586294 547274 586350
rect 547342 586294 547398 586350
rect 546970 586170 547026 586226
rect 547094 586170 547150 586226
rect 547218 586170 547274 586226
rect 547342 586170 547398 586226
rect 546970 586046 547026 586102
rect 547094 586046 547150 586102
rect 547218 586046 547274 586102
rect 547342 586046 547398 586102
rect 546970 585922 547026 585978
rect 547094 585922 547150 585978
rect 547218 585922 547274 585978
rect 547342 585922 547398 585978
rect 546970 568294 547026 568350
rect 547094 568294 547150 568350
rect 547218 568294 547274 568350
rect 547342 568294 547398 568350
rect 546970 568170 547026 568226
rect 547094 568170 547150 568226
rect 547218 568170 547274 568226
rect 547342 568170 547398 568226
rect 546970 568046 547026 568102
rect 547094 568046 547150 568102
rect 547218 568046 547274 568102
rect 547342 568046 547398 568102
rect 546970 567922 547026 567978
rect 547094 567922 547150 567978
rect 547218 567922 547274 567978
rect 547342 567922 547398 567978
rect 546970 550294 547026 550350
rect 547094 550294 547150 550350
rect 547218 550294 547274 550350
rect 547342 550294 547398 550350
rect 546970 550170 547026 550226
rect 547094 550170 547150 550226
rect 547218 550170 547274 550226
rect 547342 550170 547398 550226
rect 546970 550046 547026 550102
rect 547094 550046 547150 550102
rect 547218 550046 547274 550102
rect 547342 550046 547398 550102
rect 546970 549922 547026 549978
rect 547094 549922 547150 549978
rect 547218 549922 547274 549978
rect 547342 549922 547398 549978
rect 546970 532294 547026 532350
rect 547094 532294 547150 532350
rect 547218 532294 547274 532350
rect 547342 532294 547398 532350
rect 546970 532170 547026 532226
rect 547094 532170 547150 532226
rect 547218 532170 547274 532226
rect 547342 532170 547398 532226
rect 546970 532046 547026 532102
rect 547094 532046 547150 532102
rect 547218 532046 547274 532102
rect 547342 532046 547398 532102
rect 546970 531922 547026 531978
rect 547094 531922 547150 531978
rect 547218 531922 547274 531978
rect 547342 531922 547398 531978
rect 546970 514294 547026 514350
rect 547094 514294 547150 514350
rect 547218 514294 547274 514350
rect 547342 514294 547398 514350
rect 546970 514170 547026 514226
rect 547094 514170 547150 514226
rect 547218 514170 547274 514226
rect 547342 514170 547398 514226
rect 546970 514046 547026 514102
rect 547094 514046 547150 514102
rect 547218 514046 547274 514102
rect 547342 514046 547398 514102
rect 546970 513922 547026 513978
rect 547094 513922 547150 513978
rect 547218 513922 547274 513978
rect 547342 513922 547398 513978
rect 546970 496294 547026 496350
rect 547094 496294 547150 496350
rect 547218 496294 547274 496350
rect 547342 496294 547398 496350
rect 546970 496170 547026 496226
rect 547094 496170 547150 496226
rect 547218 496170 547274 496226
rect 547342 496170 547398 496226
rect 546970 496046 547026 496102
rect 547094 496046 547150 496102
rect 547218 496046 547274 496102
rect 547342 496046 547398 496102
rect 546970 495922 547026 495978
rect 547094 495922 547150 495978
rect 547218 495922 547274 495978
rect 547342 495922 547398 495978
rect 546970 478294 547026 478350
rect 547094 478294 547150 478350
rect 547218 478294 547274 478350
rect 547342 478294 547398 478350
rect 546970 478170 547026 478226
rect 547094 478170 547150 478226
rect 547218 478170 547274 478226
rect 547342 478170 547398 478226
rect 546970 478046 547026 478102
rect 547094 478046 547150 478102
rect 547218 478046 547274 478102
rect 547342 478046 547398 478102
rect 546970 477922 547026 477978
rect 547094 477922 547150 477978
rect 547218 477922 547274 477978
rect 547342 477922 547398 477978
rect 546970 460294 547026 460350
rect 547094 460294 547150 460350
rect 547218 460294 547274 460350
rect 547342 460294 547398 460350
rect 546970 460170 547026 460226
rect 547094 460170 547150 460226
rect 547218 460170 547274 460226
rect 547342 460170 547398 460226
rect 546970 460046 547026 460102
rect 547094 460046 547150 460102
rect 547218 460046 547274 460102
rect 547342 460046 547398 460102
rect 546970 459922 547026 459978
rect 547094 459922 547150 459978
rect 547218 459922 547274 459978
rect 547342 459922 547398 459978
rect 546970 442294 547026 442350
rect 547094 442294 547150 442350
rect 547218 442294 547274 442350
rect 547342 442294 547398 442350
rect 546970 442170 547026 442226
rect 547094 442170 547150 442226
rect 547218 442170 547274 442226
rect 547342 442170 547398 442226
rect 546970 442046 547026 442102
rect 547094 442046 547150 442102
rect 547218 442046 547274 442102
rect 547342 442046 547398 442102
rect 546970 441922 547026 441978
rect 547094 441922 547150 441978
rect 547218 441922 547274 441978
rect 547342 441922 547398 441978
rect 546970 424294 547026 424350
rect 547094 424294 547150 424350
rect 547218 424294 547274 424350
rect 547342 424294 547398 424350
rect 546970 424170 547026 424226
rect 547094 424170 547150 424226
rect 547218 424170 547274 424226
rect 547342 424170 547398 424226
rect 546970 424046 547026 424102
rect 547094 424046 547150 424102
rect 547218 424046 547274 424102
rect 547342 424046 547398 424102
rect 546970 423922 547026 423978
rect 547094 423922 547150 423978
rect 547218 423922 547274 423978
rect 547342 423922 547398 423978
rect 546970 406294 547026 406350
rect 547094 406294 547150 406350
rect 547218 406294 547274 406350
rect 547342 406294 547398 406350
rect 546970 406170 547026 406226
rect 547094 406170 547150 406226
rect 547218 406170 547274 406226
rect 547342 406170 547398 406226
rect 546970 406046 547026 406102
rect 547094 406046 547150 406102
rect 547218 406046 547274 406102
rect 547342 406046 547398 406102
rect 546970 405922 547026 405978
rect 547094 405922 547150 405978
rect 547218 405922 547274 405978
rect 547342 405922 547398 405978
rect 546970 388294 547026 388350
rect 547094 388294 547150 388350
rect 547218 388294 547274 388350
rect 547342 388294 547398 388350
rect 546970 388170 547026 388226
rect 547094 388170 547150 388226
rect 547218 388170 547274 388226
rect 547342 388170 547398 388226
rect 546970 388046 547026 388102
rect 547094 388046 547150 388102
rect 547218 388046 547274 388102
rect 547342 388046 547398 388102
rect 546970 387922 547026 387978
rect 547094 387922 547150 387978
rect 547218 387922 547274 387978
rect 547342 387922 547398 387978
rect 546970 370294 547026 370350
rect 547094 370294 547150 370350
rect 547218 370294 547274 370350
rect 547342 370294 547398 370350
rect 546970 370170 547026 370226
rect 547094 370170 547150 370226
rect 547218 370170 547274 370226
rect 547342 370170 547398 370226
rect 546970 370046 547026 370102
rect 547094 370046 547150 370102
rect 547218 370046 547274 370102
rect 547342 370046 547398 370102
rect 546970 369922 547026 369978
rect 547094 369922 547150 369978
rect 547218 369922 547274 369978
rect 547342 369922 547398 369978
rect 546970 352294 547026 352350
rect 547094 352294 547150 352350
rect 547218 352294 547274 352350
rect 547342 352294 547398 352350
rect 546970 352170 547026 352226
rect 547094 352170 547150 352226
rect 547218 352170 547274 352226
rect 547342 352170 547398 352226
rect 546970 352046 547026 352102
rect 547094 352046 547150 352102
rect 547218 352046 547274 352102
rect 547342 352046 547398 352102
rect 546970 351922 547026 351978
rect 547094 351922 547150 351978
rect 547218 351922 547274 351978
rect 547342 351922 547398 351978
rect 546970 334294 547026 334350
rect 547094 334294 547150 334350
rect 547218 334294 547274 334350
rect 547342 334294 547398 334350
rect 546970 334170 547026 334226
rect 547094 334170 547150 334226
rect 547218 334170 547274 334226
rect 547342 334170 547398 334226
rect 546970 334046 547026 334102
rect 547094 334046 547150 334102
rect 547218 334046 547274 334102
rect 547342 334046 547398 334102
rect 546970 333922 547026 333978
rect 547094 333922 547150 333978
rect 547218 333922 547274 333978
rect 547342 333922 547398 333978
rect 546970 316294 547026 316350
rect 547094 316294 547150 316350
rect 547218 316294 547274 316350
rect 547342 316294 547398 316350
rect 546970 316170 547026 316226
rect 547094 316170 547150 316226
rect 547218 316170 547274 316226
rect 547342 316170 547398 316226
rect 546970 316046 547026 316102
rect 547094 316046 547150 316102
rect 547218 316046 547274 316102
rect 547342 316046 547398 316102
rect 546970 315922 547026 315978
rect 547094 315922 547150 315978
rect 547218 315922 547274 315978
rect 547342 315922 547398 315978
rect 546970 298294 547026 298350
rect 547094 298294 547150 298350
rect 547218 298294 547274 298350
rect 547342 298294 547398 298350
rect 546970 298170 547026 298226
rect 547094 298170 547150 298226
rect 547218 298170 547274 298226
rect 547342 298170 547398 298226
rect 546970 298046 547026 298102
rect 547094 298046 547150 298102
rect 547218 298046 547274 298102
rect 547342 298046 547398 298102
rect 546970 297922 547026 297978
rect 547094 297922 547150 297978
rect 547218 297922 547274 297978
rect 547342 297922 547398 297978
rect 546970 280294 547026 280350
rect 547094 280294 547150 280350
rect 547218 280294 547274 280350
rect 547342 280294 547398 280350
rect 546970 280170 547026 280226
rect 547094 280170 547150 280226
rect 547218 280170 547274 280226
rect 547342 280170 547398 280226
rect 546970 280046 547026 280102
rect 547094 280046 547150 280102
rect 547218 280046 547274 280102
rect 547342 280046 547398 280102
rect 546970 279922 547026 279978
rect 547094 279922 547150 279978
rect 547218 279922 547274 279978
rect 547342 279922 547398 279978
rect 546970 262294 547026 262350
rect 547094 262294 547150 262350
rect 547218 262294 547274 262350
rect 547342 262294 547398 262350
rect 546970 262170 547026 262226
rect 547094 262170 547150 262226
rect 547218 262170 547274 262226
rect 547342 262170 547398 262226
rect 546970 262046 547026 262102
rect 547094 262046 547150 262102
rect 547218 262046 547274 262102
rect 547342 262046 547398 262102
rect 546970 261922 547026 261978
rect 547094 261922 547150 261978
rect 547218 261922 547274 261978
rect 547342 261922 547398 261978
rect 546970 244294 547026 244350
rect 547094 244294 547150 244350
rect 547218 244294 547274 244350
rect 547342 244294 547398 244350
rect 546970 244170 547026 244226
rect 547094 244170 547150 244226
rect 547218 244170 547274 244226
rect 547342 244170 547398 244226
rect 546970 244046 547026 244102
rect 547094 244046 547150 244102
rect 547218 244046 547274 244102
rect 547342 244046 547398 244102
rect 546970 243922 547026 243978
rect 547094 243922 547150 243978
rect 547218 243922 547274 243978
rect 547342 243922 547398 243978
rect 546970 226294 547026 226350
rect 547094 226294 547150 226350
rect 547218 226294 547274 226350
rect 547342 226294 547398 226350
rect 546970 226170 547026 226226
rect 547094 226170 547150 226226
rect 547218 226170 547274 226226
rect 547342 226170 547398 226226
rect 546970 226046 547026 226102
rect 547094 226046 547150 226102
rect 547218 226046 547274 226102
rect 547342 226046 547398 226102
rect 546970 225922 547026 225978
rect 547094 225922 547150 225978
rect 547218 225922 547274 225978
rect 547342 225922 547398 225978
rect 546970 208294 547026 208350
rect 547094 208294 547150 208350
rect 547218 208294 547274 208350
rect 547342 208294 547398 208350
rect 546970 208170 547026 208226
rect 547094 208170 547150 208226
rect 547218 208170 547274 208226
rect 547342 208170 547398 208226
rect 546970 208046 547026 208102
rect 547094 208046 547150 208102
rect 547218 208046 547274 208102
rect 547342 208046 547398 208102
rect 546970 207922 547026 207978
rect 547094 207922 547150 207978
rect 547218 207922 547274 207978
rect 547342 207922 547398 207978
rect 546970 190294 547026 190350
rect 547094 190294 547150 190350
rect 547218 190294 547274 190350
rect 547342 190294 547398 190350
rect 546970 190170 547026 190226
rect 547094 190170 547150 190226
rect 547218 190170 547274 190226
rect 547342 190170 547398 190226
rect 546970 190046 547026 190102
rect 547094 190046 547150 190102
rect 547218 190046 547274 190102
rect 547342 190046 547398 190102
rect 546970 189922 547026 189978
rect 547094 189922 547150 189978
rect 547218 189922 547274 189978
rect 547342 189922 547398 189978
rect 546970 172294 547026 172350
rect 547094 172294 547150 172350
rect 547218 172294 547274 172350
rect 547342 172294 547398 172350
rect 546970 172170 547026 172226
rect 547094 172170 547150 172226
rect 547218 172170 547274 172226
rect 547342 172170 547398 172226
rect 546970 172046 547026 172102
rect 547094 172046 547150 172102
rect 547218 172046 547274 172102
rect 547342 172046 547398 172102
rect 546970 171922 547026 171978
rect 547094 171922 547150 171978
rect 547218 171922 547274 171978
rect 547342 171922 547398 171978
rect 546970 154294 547026 154350
rect 547094 154294 547150 154350
rect 547218 154294 547274 154350
rect 547342 154294 547398 154350
rect 546970 154170 547026 154226
rect 547094 154170 547150 154226
rect 547218 154170 547274 154226
rect 547342 154170 547398 154226
rect 546970 154046 547026 154102
rect 547094 154046 547150 154102
rect 547218 154046 547274 154102
rect 547342 154046 547398 154102
rect 546970 153922 547026 153978
rect 547094 153922 547150 153978
rect 547218 153922 547274 153978
rect 547342 153922 547398 153978
rect 546970 136294 547026 136350
rect 547094 136294 547150 136350
rect 547218 136294 547274 136350
rect 547342 136294 547398 136350
rect 546970 136170 547026 136226
rect 547094 136170 547150 136226
rect 547218 136170 547274 136226
rect 547342 136170 547398 136226
rect 546970 136046 547026 136102
rect 547094 136046 547150 136102
rect 547218 136046 547274 136102
rect 547342 136046 547398 136102
rect 546970 135922 547026 135978
rect 547094 135922 547150 135978
rect 547218 135922 547274 135978
rect 547342 135922 547398 135978
rect 546970 118294 547026 118350
rect 547094 118294 547150 118350
rect 547218 118294 547274 118350
rect 547342 118294 547398 118350
rect 546970 118170 547026 118226
rect 547094 118170 547150 118226
rect 547218 118170 547274 118226
rect 547342 118170 547398 118226
rect 546970 118046 547026 118102
rect 547094 118046 547150 118102
rect 547218 118046 547274 118102
rect 547342 118046 547398 118102
rect 546970 117922 547026 117978
rect 547094 117922 547150 117978
rect 547218 117922 547274 117978
rect 547342 117922 547398 117978
rect 546970 100294 547026 100350
rect 547094 100294 547150 100350
rect 547218 100294 547274 100350
rect 547342 100294 547398 100350
rect 546970 100170 547026 100226
rect 547094 100170 547150 100226
rect 547218 100170 547274 100226
rect 547342 100170 547398 100226
rect 546970 100046 547026 100102
rect 547094 100046 547150 100102
rect 547218 100046 547274 100102
rect 547342 100046 547398 100102
rect 546970 99922 547026 99978
rect 547094 99922 547150 99978
rect 547218 99922 547274 99978
rect 547342 99922 547398 99978
rect 546970 82294 547026 82350
rect 547094 82294 547150 82350
rect 547218 82294 547274 82350
rect 547342 82294 547398 82350
rect 546970 82170 547026 82226
rect 547094 82170 547150 82226
rect 547218 82170 547274 82226
rect 547342 82170 547398 82226
rect 546970 82046 547026 82102
rect 547094 82046 547150 82102
rect 547218 82046 547274 82102
rect 547342 82046 547398 82102
rect 546970 81922 547026 81978
rect 547094 81922 547150 81978
rect 547218 81922 547274 81978
rect 547342 81922 547398 81978
rect 546970 64294 547026 64350
rect 547094 64294 547150 64350
rect 547218 64294 547274 64350
rect 547342 64294 547398 64350
rect 546970 64170 547026 64226
rect 547094 64170 547150 64226
rect 547218 64170 547274 64226
rect 547342 64170 547398 64226
rect 546970 64046 547026 64102
rect 547094 64046 547150 64102
rect 547218 64046 547274 64102
rect 547342 64046 547398 64102
rect 546970 63922 547026 63978
rect 547094 63922 547150 63978
rect 547218 63922 547274 63978
rect 547342 63922 547398 63978
rect 546970 46294 547026 46350
rect 547094 46294 547150 46350
rect 547218 46294 547274 46350
rect 547342 46294 547398 46350
rect 546970 46170 547026 46226
rect 547094 46170 547150 46226
rect 547218 46170 547274 46226
rect 547342 46170 547398 46226
rect 546970 46046 547026 46102
rect 547094 46046 547150 46102
rect 547218 46046 547274 46102
rect 547342 46046 547398 46102
rect 546970 45922 547026 45978
rect 547094 45922 547150 45978
rect 547218 45922 547274 45978
rect 547342 45922 547398 45978
rect 546970 28294 547026 28350
rect 547094 28294 547150 28350
rect 547218 28294 547274 28350
rect 547342 28294 547398 28350
rect 546970 28170 547026 28226
rect 547094 28170 547150 28226
rect 547218 28170 547274 28226
rect 547342 28170 547398 28226
rect 546970 28046 547026 28102
rect 547094 28046 547150 28102
rect 547218 28046 547274 28102
rect 547342 28046 547398 28102
rect 546970 27922 547026 27978
rect 547094 27922 547150 27978
rect 547218 27922 547274 27978
rect 547342 27922 547398 27978
rect 546970 10294 547026 10350
rect 547094 10294 547150 10350
rect 547218 10294 547274 10350
rect 547342 10294 547398 10350
rect 546970 10170 547026 10226
rect 547094 10170 547150 10226
rect 547218 10170 547274 10226
rect 547342 10170 547398 10226
rect 546970 10046 547026 10102
rect 547094 10046 547150 10102
rect 547218 10046 547274 10102
rect 547342 10046 547398 10102
rect 546970 9922 547026 9978
rect 547094 9922 547150 9978
rect 547218 9922 547274 9978
rect 547342 9922 547398 9978
rect 546970 -1176 547026 -1120
rect 547094 -1176 547150 -1120
rect 547218 -1176 547274 -1120
rect 547342 -1176 547398 -1120
rect 546970 -1300 547026 -1244
rect 547094 -1300 547150 -1244
rect 547218 -1300 547274 -1244
rect 547342 -1300 547398 -1244
rect 546970 -1424 547026 -1368
rect 547094 -1424 547150 -1368
rect 547218 -1424 547274 -1368
rect 547342 -1424 547398 -1368
rect 546970 -1548 547026 -1492
rect 547094 -1548 547150 -1492
rect 547218 -1548 547274 -1492
rect 547342 -1548 547398 -1492
rect 561250 597156 561306 597212
rect 561374 597156 561430 597212
rect 561498 597156 561554 597212
rect 561622 597156 561678 597212
rect 561250 597032 561306 597088
rect 561374 597032 561430 597088
rect 561498 597032 561554 597088
rect 561622 597032 561678 597088
rect 561250 596908 561306 596964
rect 561374 596908 561430 596964
rect 561498 596908 561554 596964
rect 561622 596908 561678 596964
rect 561250 596784 561306 596840
rect 561374 596784 561430 596840
rect 561498 596784 561554 596840
rect 561622 596784 561678 596840
rect 561250 580294 561306 580350
rect 561374 580294 561430 580350
rect 561498 580294 561554 580350
rect 561622 580294 561678 580350
rect 561250 580170 561306 580226
rect 561374 580170 561430 580226
rect 561498 580170 561554 580226
rect 561622 580170 561678 580226
rect 561250 580046 561306 580102
rect 561374 580046 561430 580102
rect 561498 580046 561554 580102
rect 561622 580046 561678 580102
rect 561250 579922 561306 579978
rect 561374 579922 561430 579978
rect 561498 579922 561554 579978
rect 561622 579922 561678 579978
rect 561250 562294 561306 562350
rect 561374 562294 561430 562350
rect 561498 562294 561554 562350
rect 561622 562294 561678 562350
rect 561250 562170 561306 562226
rect 561374 562170 561430 562226
rect 561498 562170 561554 562226
rect 561622 562170 561678 562226
rect 561250 562046 561306 562102
rect 561374 562046 561430 562102
rect 561498 562046 561554 562102
rect 561622 562046 561678 562102
rect 561250 561922 561306 561978
rect 561374 561922 561430 561978
rect 561498 561922 561554 561978
rect 561622 561922 561678 561978
rect 561250 544294 561306 544350
rect 561374 544294 561430 544350
rect 561498 544294 561554 544350
rect 561622 544294 561678 544350
rect 561250 544170 561306 544226
rect 561374 544170 561430 544226
rect 561498 544170 561554 544226
rect 561622 544170 561678 544226
rect 561250 544046 561306 544102
rect 561374 544046 561430 544102
rect 561498 544046 561554 544102
rect 561622 544046 561678 544102
rect 561250 543922 561306 543978
rect 561374 543922 561430 543978
rect 561498 543922 561554 543978
rect 561622 543922 561678 543978
rect 561250 526294 561306 526350
rect 561374 526294 561430 526350
rect 561498 526294 561554 526350
rect 561622 526294 561678 526350
rect 561250 526170 561306 526226
rect 561374 526170 561430 526226
rect 561498 526170 561554 526226
rect 561622 526170 561678 526226
rect 561250 526046 561306 526102
rect 561374 526046 561430 526102
rect 561498 526046 561554 526102
rect 561622 526046 561678 526102
rect 561250 525922 561306 525978
rect 561374 525922 561430 525978
rect 561498 525922 561554 525978
rect 561622 525922 561678 525978
rect 561250 508294 561306 508350
rect 561374 508294 561430 508350
rect 561498 508294 561554 508350
rect 561622 508294 561678 508350
rect 561250 508170 561306 508226
rect 561374 508170 561430 508226
rect 561498 508170 561554 508226
rect 561622 508170 561678 508226
rect 561250 508046 561306 508102
rect 561374 508046 561430 508102
rect 561498 508046 561554 508102
rect 561622 508046 561678 508102
rect 561250 507922 561306 507978
rect 561374 507922 561430 507978
rect 561498 507922 561554 507978
rect 561622 507922 561678 507978
rect 561250 490294 561306 490350
rect 561374 490294 561430 490350
rect 561498 490294 561554 490350
rect 561622 490294 561678 490350
rect 561250 490170 561306 490226
rect 561374 490170 561430 490226
rect 561498 490170 561554 490226
rect 561622 490170 561678 490226
rect 561250 490046 561306 490102
rect 561374 490046 561430 490102
rect 561498 490046 561554 490102
rect 561622 490046 561678 490102
rect 561250 489922 561306 489978
rect 561374 489922 561430 489978
rect 561498 489922 561554 489978
rect 561622 489922 561678 489978
rect 561250 472294 561306 472350
rect 561374 472294 561430 472350
rect 561498 472294 561554 472350
rect 561622 472294 561678 472350
rect 561250 472170 561306 472226
rect 561374 472170 561430 472226
rect 561498 472170 561554 472226
rect 561622 472170 561678 472226
rect 561250 472046 561306 472102
rect 561374 472046 561430 472102
rect 561498 472046 561554 472102
rect 561622 472046 561678 472102
rect 561250 471922 561306 471978
rect 561374 471922 561430 471978
rect 561498 471922 561554 471978
rect 561622 471922 561678 471978
rect 561250 454294 561306 454350
rect 561374 454294 561430 454350
rect 561498 454294 561554 454350
rect 561622 454294 561678 454350
rect 561250 454170 561306 454226
rect 561374 454170 561430 454226
rect 561498 454170 561554 454226
rect 561622 454170 561678 454226
rect 561250 454046 561306 454102
rect 561374 454046 561430 454102
rect 561498 454046 561554 454102
rect 561622 454046 561678 454102
rect 561250 453922 561306 453978
rect 561374 453922 561430 453978
rect 561498 453922 561554 453978
rect 561622 453922 561678 453978
rect 561250 436294 561306 436350
rect 561374 436294 561430 436350
rect 561498 436294 561554 436350
rect 561622 436294 561678 436350
rect 561250 436170 561306 436226
rect 561374 436170 561430 436226
rect 561498 436170 561554 436226
rect 561622 436170 561678 436226
rect 561250 436046 561306 436102
rect 561374 436046 561430 436102
rect 561498 436046 561554 436102
rect 561622 436046 561678 436102
rect 561250 435922 561306 435978
rect 561374 435922 561430 435978
rect 561498 435922 561554 435978
rect 561622 435922 561678 435978
rect 561250 418294 561306 418350
rect 561374 418294 561430 418350
rect 561498 418294 561554 418350
rect 561622 418294 561678 418350
rect 561250 418170 561306 418226
rect 561374 418170 561430 418226
rect 561498 418170 561554 418226
rect 561622 418170 561678 418226
rect 561250 418046 561306 418102
rect 561374 418046 561430 418102
rect 561498 418046 561554 418102
rect 561622 418046 561678 418102
rect 561250 417922 561306 417978
rect 561374 417922 561430 417978
rect 561498 417922 561554 417978
rect 561622 417922 561678 417978
rect 561250 400294 561306 400350
rect 561374 400294 561430 400350
rect 561498 400294 561554 400350
rect 561622 400294 561678 400350
rect 561250 400170 561306 400226
rect 561374 400170 561430 400226
rect 561498 400170 561554 400226
rect 561622 400170 561678 400226
rect 561250 400046 561306 400102
rect 561374 400046 561430 400102
rect 561498 400046 561554 400102
rect 561622 400046 561678 400102
rect 561250 399922 561306 399978
rect 561374 399922 561430 399978
rect 561498 399922 561554 399978
rect 561622 399922 561678 399978
rect 561250 382294 561306 382350
rect 561374 382294 561430 382350
rect 561498 382294 561554 382350
rect 561622 382294 561678 382350
rect 561250 382170 561306 382226
rect 561374 382170 561430 382226
rect 561498 382170 561554 382226
rect 561622 382170 561678 382226
rect 561250 382046 561306 382102
rect 561374 382046 561430 382102
rect 561498 382046 561554 382102
rect 561622 382046 561678 382102
rect 561250 381922 561306 381978
rect 561374 381922 561430 381978
rect 561498 381922 561554 381978
rect 561622 381922 561678 381978
rect 561250 364294 561306 364350
rect 561374 364294 561430 364350
rect 561498 364294 561554 364350
rect 561622 364294 561678 364350
rect 561250 364170 561306 364226
rect 561374 364170 561430 364226
rect 561498 364170 561554 364226
rect 561622 364170 561678 364226
rect 561250 364046 561306 364102
rect 561374 364046 561430 364102
rect 561498 364046 561554 364102
rect 561622 364046 561678 364102
rect 561250 363922 561306 363978
rect 561374 363922 561430 363978
rect 561498 363922 561554 363978
rect 561622 363922 561678 363978
rect 561250 346294 561306 346350
rect 561374 346294 561430 346350
rect 561498 346294 561554 346350
rect 561622 346294 561678 346350
rect 561250 346170 561306 346226
rect 561374 346170 561430 346226
rect 561498 346170 561554 346226
rect 561622 346170 561678 346226
rect 561250 346046 561306 346102
rect 561374 346046 561430 346102
rect 561498 346046 561554 346102
rect 561622 346046 561678 346102
rect 561250 345922 561306 345978
rect 561374 345922 561430 345978
rect 561498 345922 561554 345978
rect 561622 345922 561678 345978
rect 561250 328294 561306 328350
rect 561374 328294 561430 328350
rect 561498 328294 561554 328350
rect 561622 328294 561678 328350
rect 561250 328170 561306 328226
rect 561374 328170 561430 328226
rect 561498 328170 561554 328226
rect 561622 328170 561678 328226
rect 561250 328046 561306 328102
rect 561374 328046 561430 328102
rect 561498 328046 561554 328102
rect 561622 328046 561678 328102
rect 561250 327922 561306 327978
rect 561374 327922 561430 327978
rect 561498 327922 561554 327978
rect 561622 327922 561678 327978
rect 561250 310294 561306 310350
rect 561374 310294 561430 310350
rect 561498 310294 561554 310350
rect 561622 310294 561678 310350
rect 561250 310170 561306 310226
rect 561374 310170 561430 310226
rect 561498 310170 561554 310226
rect 561622 310170 561678 310226
rect 561250 310046 561306 310102
rect 561374 310046 561430 310102
rect 561498 310046 561554 310102
rect 561622 310046 561678 310102
rect 561250 309922 561306 309978
rect 561374 309922 561430 309978
rect 561498 309922 561554 309978
rect 561622 309922 561678 309978
rect 561250 292294 561306 292350
rect 561374 292294 561430 292350
rect 561498 292294 561554 292350
rect 561622 292294 561678 292350
rect 561250 292170 561306 292226
rect 561374 292170 561430 292226
rect 561498 292170 561554 292226
rect 561622 292170 561678 292226
rect 561250 292046 561306 292102
rect 561374 292046 561430 292102
rect 561498 292046 561554 292102
rect 561622 292046 561678 292102
rect 561250 291922 561306 291978
rect 561374 291922 561430 291978
rect 561498 291922 561554 291978
rect 561622 291922 561678 291978
rect 561250 274294 561306 274350
rect 561374 274294 561430 274350
rect 561498 274294 561554 274350
rect 561622 274294 561678 274350
rect 561250 274170 561306 274226
rect 561374 274170 561430 274226
rect 561498 274170 561554 274226
rect 561622 274170 561678 274226
rect 561250 274046 561306 274102
rect 561374 274046 561430 274102
rect 561498 274046 561554 274102
rect 561622 274046 561678 274102
rect 561250 273922 561306 273978
rect 561374 273922 561430 273978
rect 561498 273922 561554 273978
rect 561622 273922 561678 273978
rect 561250 256294 561306 256350
rect 561374 256294 561430 256350
rect 561498 256294 561554 256350
rect 561622 256294 561678 256350
rect 561250 256170 561306 256226
rect 561374 256170 561430 256226
rect 561498 256170 561554 256226
rect 561622 256170 561678 256226
rect 561250 256046 561306 256102
rect 561374 256046 561430 256102
rect 561498 256046 561554 256102
rect 561622 256046 561678 256102
rect 561250 255922 561306 255978
rect 561374 255922 561430 255978
rect 561498 255922 561554 255978
rect 561622 255922 561678 255978
rect 561250 238294 561306 238350
rect 561374 238294 561430 238350
rect 561498 238294 561554 238350
rect 561622 238294 561678 238350
rect 561250 238170 561306 238226
rect 561374 238170 561430 238226
rect 561498 238170 561554 238226
rect 561622 238170 561678 238226
rect 561250 238046 561306 238102
rect 561374 238046 561430 238102
rect 561498 238046 561554 238102
rect 561622 238046 561678 238102
rect 561250 237922 561306 237978
rect 561374 237922 561430 237978
rect 561498 237922 561554 237978
rect 561622 237922 561678 237978
rect 561250 220294 561306 220350
rect 561374 220294 561430 220350
rect 561498 220294 561554 220350
rect 561622 220294 561678 220350
rect 561250 220170 561306 220226
rect 561374 220170 561430 220226
rect 561498 220170 561554 220226
rect 561622 220170 561678 220226
rect 561250 220046 561306 220102
rect 561374 220046 561430 220102
rect 561498 220046 561554 220102
rect 561622 220046 561678 220102
rect 561250 219922 561306 219978
rect 561374 219922 561430 219978
rect 561498 219922 561554 219978
rect 561622 219922 561678 219978
rect 561250 202294 561306 202350
rect 561374 202294 561430 202350
rect 561498 202294 561554 202350
rect 561622 202294 561678 202350
rect 561250 202170 561306 202226
rect 561374 202170 561430 202226
rect 561498 202170 561554 202226
rect 561622 202170 561678 202226
rect 561250 202046 561306 202102
rect 561374 202046 561430 202102
rect 561498 202046 561554 202102
rect 561622 202046 561678 202102
rect 561250 201922 561306 201978
rect 561374 201922 561430 201978
rect 561498 201922 561554 201978
rect 561622 201922 561678 201978
rect 561250 184294 561306 184350
rect 561374 184294 561430 184350
rect 561498 184294 561554 184350
rect 561622 184294 561678 184350
rect 561250 184170 561306 184226
rect 561374 184170 561430 184226
rect 561498 184170 561554 184226
rect 561622 184170 561678 184226
rect 561250 184046 561306 184102
rect 561374 184046 561430 184102
rect 561498 184046 561554 184102
rect 561622 184046 561678 184102
rect 561250 183922 561306 183978
rect 561374 183922 561430 183978
rect 561498 183922 561554 183978
rect 561622 183922 561678 183978
rect 561250 166294 561306 166350
rect 561374 166294 561430 166350
rect 561498 166294 561554 166350
rect 561622 166294 561678 166350
rect 561250 166170 561306 166226
rect 561374 166170 561430 166226
rect 561498 166170 561554 166226
rect 561622 166170 561678 166226
rect 561250 166046 561306 166102
rect 561374 166046 561430 166102
rect 561498 166046 561554 166102
rect 561622 166046 561678 166102
rect 561250 165922 561306 165978
rect 561374 165922 561430 165978
rect 561498 165922 561554 165978
rect 561622 165922 561678 165978
rect 561250 148294 561306 148350
rect 561374 148294 561430 148350
rect 561498 148294 561554 148350
rect 561622 148294 561678 148350
rect 561250 148170 561306 148226
rect 561374 148170 561430 148226
rect 561498 148170 561554 148226
rect 561622 148170 561678 148226
rect 561250 148046 561306 148102
rect 561374 148046 561430 148102
rect 561498 148046 561554 148102
rect 561622 148046 561678 148102
rect 561250 147922 561306 147978
rect 561374 147922 561430 147978
rect 561498 147922 561554 147978
rect 561622 147922 561678 147978
rect 561250 130294 561306 130350
rect 561374 130294 561430 130350
rect 561498 130294 561554 130350
rect 561622 130294 561678 130350
rect 561250 130170 561306 130226
rect 561374 130170 561430 130226
rect 561498 130170 561554 130226
rect 561622 130170 561678 130226
rect 561250 130046 561306 130102
rect 561374 130046 561430 130102
rect 561498 130046 561554 130102
rect 561622 130046 561678 130102
rect 561250 129922 561306 129978
rect 561374 129922 561430 129978
rect 561498 129922 561554 129978
rect 561622 129922 561678 129978
rect 561250 112294 561306 112350
rect 561374 112294 561430 112350
rect 561498 112294 561554 112350
rect 561622 112294 561678 112350
rect 561250 112170 561306 112226
rect 561374 112170 561430 112226
rect 561498 112170 561554 112226
rect 561622 112170 561678 112226
rect 561250 112046 561306 112102
rect 561374 112046 561430 112102
rect 561498 112046 561554 112102
rect 561622 112046 561678 112102
rect 561250 111922 561306 111978
rect 561374 111922 561430 111978
rect 561498 111922 561554 111978
rect 561622 111922 561678 111978
rect 561250 94294 561306 94350
rect 561374 94294 561430 94350
rect 561498 94294 561554 94350
rect 561622 94294 561678 94350
rect 561250 94170 561306 94226
rect 561374 94170 561430 94226
rect 561498 94170 561554 94226
rect 561622 94170 561678 94226
rect 561250 94046 561306 94102
rect 561374 94046 561430 94102
rect 561498 94046 561554 94102
rect 561622 94046 561678 94102
rect 561250 93922 561306 93978
rect 561374 93922 561430 93978
rect 561498 93922 561554 93978
rect 561622 93922 561678 93978
rect 561250 76294 561306 76350
rect 561374 76294 561430 76350
rect 561498 76294 561554 76350
rect 561622 76294 561678 76350
rect 561250 76170 561306 76226
rect 561374 76170 561430 76226
rect 561498 76170 561554 76226
rect 561622 76170 561678 76226
rect 561250 76046 561306 76102
rect 561374 76046 561430 76102
rect 561498 76046 561554 76102
rect 561622 76046 561678 76102
rect 561250 75922 561306 75978
rect 561374 75922 561430 75978
rect 561498 75922 561554 75978
rect 561622 75922 561678 75978
rect 561250 58294 561306 58350
rect 561374 58294 561430 58350
rect 561498 58294 561554 58350
rect 561622 58294 561678 58350
rect 561250 58170 561306 58226
rect 561374 58170 561430 58226
rect 561498 58170 561554 58226
rect 561622 58170 561678 58226
rect 561250 58046 561306 58102
rect 561374 58046 561430 58102
rect 561498 58046 561554 58102
rect 561622 58046 561678 58102
rect 561250 57922 561306 57978
rect 561374 57922 561430 57978
rect 561498 57922 561554 57978
rect 561622 57922 561678 57978
rect 561250 40294 561306 40350
rect 561374 40294 561430 40350
rect 561498 40294 561554 40350
rect 561622 40294 561678 40350
rect 561250 40170 561306 40226
rect 561374 40170 561430 40226
rect 561498 40170 561554 40226
rect 561622 40170 561678 40226
rect 561250 40046 561306 40102
rect 561374 40046 561430 40102
rect 561498 40046 561554 40102
rect 561622 40046 561678 40102
rect 561250 39922 561306 39978
rect 561374 39922 561430 39978
rect 561498 39922 561554 39978
rect 561622 39922 561678 39978
rect 561250 22294 561306 22350
rect 561374 22294 561430 22350
rect 561498 22294 561554 22350
rect 561622 22294 561678 22350
rect 561250 22170 561306 22226
rect 561374 22170 561430 22226
rect 561498 22170 561554 22226
rect 561622 22170 561678 22226
rect 561250 22046 561306 22102
rect 561374 22046 561430 22102
rect 561498 22046 561554 22102
rect 561622 22046 561678 22102
rect 561250 21922 561306 21978
rect 561374 21922 561430 21978
rect 561498 21922 561554 21978
rect 561622 21922 561678 21978
rect 561250 4294 561306 4350
rect 561374 4294 561430 4350
rect 561498 4294 561554 4350
rect 561622 4294 561678 4350
rect 561250 4170 561306 4226
rect 561374 4170 561430 4226
rect 561498 4170 561554 4226
rect 561622 4170 561678 4226
rect 561250 4046 561306 4102
rect 561374 4046 561430 4102
rect 561498 4046 561554 4102
rect 561622 4046 561678 4102
rect 561250 3922 561306 3978
rect 561374 3922 561430 3978
rect 561498 3922 561554 3978
rect 561622 3922 561678 3978
rect 561250 -216 561306 -160
rect 561374 -216 561430 -160
rect 561498 -216 561554 -160
rect 561622 -216 561678 -160
rect 561250 -340 561306 -284
rect 561374 -340 561430 -284
rect 561498 -340 561554 -284
rect 561622 -340 561678 -284
rect 561250 -464 561306 -408
rect 561374 -464 561430 -408
rect 561498 -464 561554 -408
rect 561622 -464 561678 -408
rect 561250 -588 561306 -532
rect 561374 -588 561430 -532
rect 561498 -588 561554 -532
rect 561622 -588 561678 -532
rect 564970 598116 565026 598172
rect 565094 598116 565150 598172
rect 565218 598116 565274 598172
rect 565342 598116 565398 598172
rect 564970 597992 565026 598048
rect 565094 597992 565150 598048
rect 565218 597992 565274 598048
rect 565342 597992 565398 598048
rect 564970 597868 565026 597924
rect 565094 597868 565150 597924
rect 565218 597868 565274 597924
rect 565342 597868 565398 597924
rect 564970 597744 565026 597800
rect 565094 597744 565150 597800
rect 565218 597744 565274 597800
rect 565342 597744 565398 597800
rect 564970 586294 565026 586350
rect 565094 586294 565150 586350
rect 565218 586294 565274 586350
rect 565342 586294 565398 586350
rect 564970 586170 565026 586226
rect 565094 586170 565150 586226
rect 565218 586170 565274 586226
rect 565342 586170 565398 586226
rect 564970 586046 565026 586102
rect 565094 586046 565150 586102
rect 565218 586046 565274 586102
rect 565342 586046 565398 586102
rect 564970 585922 565026 585978
rect 565094 585922 565150 585978
rect 565218 585922 565274 585978
rect 565342 585922 565398 585978
rect 564970 568294 565026 568350
rect 565094 568294 565150 568350
rect 565218 568294 565274 568350
rect 565342 568294 565398 568350
rect 564970 568170 565026 568226
rect 565094 568170 565150 568226
rect 565218 568170 565274 568226
rect 565342 568170 565398 568226
rect 564970 568046 565026 568102
rect 565094 568046 565150 568102
rect 565218 568046 565274 568102
rect 565342 568046 565398 568102
rect 564970 567922 565026 567978
rect 565094 567922 565150 567978
rect 565218 567922 565274 567978
rect 565342 567922 565398 567978
rect 564970 550294 565026 550350
rect 565094 550294 565150 550350
rect 565218 550294 565274 550350
rect 565342 550294 565398 550350
rect 564970 550170 565026 550226
rect 565094 550170 565150 550226
rect 565218 550170 565274 550226
rect 565342 550170 565398 550226
rect 564970 550046 565026 550102
rect 565094 550046 565150 550102
rect 565218 550046 565274 550102
rect 565342 550046 565398 550102
rect 564970 549922 565026 549978
rect 565094 549922 565150 549978
rect 565218 549922 565274 549978
rect 565342 549922 565398 549978
rect 564970 532294 565026 532350
rect 565094 532294 565150 532350
rect 565218 532294 565274 532350
rect 565342 532294 565398 532350
rect 564970 532170 565026 532226
rect 565094 532170 565150 532226
rect 565218 532170 565274 532226
rect 565342 532170 565398 532226
rect 564970 532046 565026 532102
rect 565094 532046 565150 532102
rect 565218 532046 565274 532102
rect 565342 532046 565398 532102
rect 564970 531922 565026 531978
rect 565094 531922 565150 531978
rect 565218 531922 565274 531978
rect 565342 531922 565398 531978
rect 564970 514294 565026 514350
rect 565094 514294 565150 514350
rect 565218 514294 565274 514350
rect 565342 514294 565398 514350
rect 564970 514170 565026 514226
rect 565094 514170 565150 514226
rect 565218 514170 565274 514226
rect 565342 514170 565398 514226
rect 564970 514046 565026 514102
rect 565094 514046 565150 514102
rect 565218 514046 565274 514102
rect 565342 514046 565398 514102
rect 564970 513922 565026 513978
rect 565094 513922 565150 513978
rect 565218 513922 565274 513978
rect 565342 513922 565398 513978
rect 564970 496294 565026 496350
rect 565094 496294 565150 496350
rect 565218 496294 565274 496350
rect 565342 496294 565398 496350
rect 564970 496170 565026 496226
rect 565094 496170 565150 496226
rect 565218 496170 565274 496226
rect 565342 496170 565398 496226
rect 564970 496046 565026 496102
rect 565094 496046 565150 496102
rect 565218 496046 565274 496102
rect 565342 496046 565398 496102
rect 564970 495922 565026 495978
rect 565094 495922 565150 495978
rect 565218 495922 565274 495978
rect 565342 495922 565398 495978
rect 564970 478294 565026 478350
rect 565094 478294 565150 478350
rect 565218 478294 565274 478350
rect 565342 478294 565398 478350
rect 564970 478170 565026 478226
rect 565094 478170 565150 478226
rect 565218 478170 565274 478226
rect 565342 478170 565398 478226
rect 564970 478046 565026 478102
rect 565094 478046 565150 478102
rect 565218 478046 565274 478102
rect 565342 478046 565398 478102
rect 564970 477922 565026 477978
rect 565094 477922 565150 477978
rect 565218 477922 565274 477978
rect 565342 477922 565398 477978
rect 564970 460294 565026 460350
rect 565094 460294 565150 460350
rect 565218 460294 565274 460350
rect 565342 460294 565398 460350
rect 564970 460170 565026 460226
rect 565094 460170 565150 460226
rect 565218 460170 565274 460226
rect 565342 460170 565398 460226
rect 564970 460046 565026 460102
rect 565094 460046 565150 460102
rect 565218 460046 565274 460102
rect 565342 460046 565398 460102
rect 564970 459922 565026 459978
rect 565094 459922 565150 459978
rect 565218 459922 565274 459978
rect 565342 459922 565398 459978
rect 564970 442294 565026 442350
rect 565094 442294 565150 442350
rect 565218 442294 565274 442350
rect 565342 442294 565398 442350
rect 564970 442170 565026 442226
rect 565094 442170 565150 442226
rect 565218 442170 565274 442226
rect 565342 442170 565398 442226
rect 564970 442046 565026 442102
rect 565094 442046 565150 442102
rect 565218 442046 565274 442102
rect 565342 442046 565398 442102
rect 564970 441922 565026 441978
rect 565094 441922 565150 441978
rect 565218 441922 565274 441978
rect 565342 441922 565398 441978
rect 564970 424294 565026 424350
rect 565094 424294 565150 424350
rect 565218 424294 565274 424350
rect 565342 424294 565398 424350
rect 564970 424170 565026 424226
rect 565094 424170 565150 424226
rect 565218 424170 565274 424226
rect 565342 424170 565398 424226
rect 564970 424046 565026 424102
rect 565094 424046 565150 424102
rect 565218 424046 565274 424102
rect 565342 424046 565398 424102
rect 564970 423922 565026 423978
rect 565094 423922 565150 423978
rect 565218 423922 565274 423978
rect 565342 423922 565398 423978
rect 564970 406294 565026 406350
rect 565094 406294 565150 406350
rect 565218 406294 565274 406350
rect 565342 406294 565398 406350
rect 564970 406170 565026 406226
rect 565094 406170 565150 406226
rect 565218 406170 565274 406226
rect 565342 406170 565398 406226
rect 564970 406046 565026 406102
rect 565094 406046 565150 406102
rect 565218 406046 565274 406102
rect 565342 406046 565398 406102
rect 564970 405922 565026 405978
rect 565094 405922 565150 405978
rect 565218 405922 565274 405978
rect 565342 405922 565398 405978
rect 564970 388294 565026 388350
rect 565094 388294 565150 388350
rect 565218 388294 565274 388350
rect 565342 388294 565398 388350
rect 564970 388170 565026 388226
rect 565094 388170 565150 388226
rect 565218 388170 565274 388226
rect 565342 388170 565398 388226
rect 564970 388046 565026 388102
rect 565094 388046 565150 388102
rect 565218 388046 565274 388102
rect 565342 388046 565398 388102
rect 564970 387922 565026 387978
rect 565094 387922 565150 387978
rect 565218 387922 565274 387978
rect 565342 387922 565398 387978
rect 564970 370294 565026 370350
rect 565094 370294 565150 370350
rect 565218 370294 565274 370350
rect 565342 370294 565398 370350
rect 564970 370170 565026 370226
rect 565094 370170 565150 370226
rect 565218 370170 565274 370226
rect 565342 370170 565398 370226
rect 564970 370046 565026 370102
rect 565094 370046 565150 370102
rect 565218 370046 565274 370102
rect 565342 370046 565398 370102
rect 564970 369922 565026 369978
rect 565094 369922 565150 369978
rect 565218 369922 565274 369978
rect 565342 369922 565398 369978
rect 564970 352294 565026 352350
rect 565094 352294 565150 352350
rect 565218 352294 565274 352350
rect 565342 352294 565398 352350
rect 564970 352170 565026 352226
rect 565094 352170 565150 352226
rect 565218 352170 565274 352226
rect 565342 352170 565398 352226
rect 564970 352046 565026 352102
rect 565094 352046 565150 352102
rect 565218 352046 565274 352102
rect 565342 352046 565398 352102
rect 564970 351922 565026 351978
rect 565094 351922 565150 351978
rect 565218 351922 565274 351978
rect 565342 351922 565398 351978
rect 564970 334294 565026 334350
rect 565094 334294 565150 334350
rect 565218 334294 565274 334350
rect 565342 334294 565398 334350
rect 564970 334170 565026 334226
rect 565094 334170 565150 334226
rect 565218 334170 565274 334226
rect 565342 334170 565398 334226
rect 564970 334046 565026 334102
rect 565094 334046 565150 334102
rect 565218 334046 565274 334102
rect 565342 334046 565398 334102
rect 564970 333922 565026 333978
rect 565094 333922 565150 333978
rect 565218 333922 565274 333978
rect 565342 333922 565398 333978
rect 564970 316294 565026 316350
rect 565094 316294 565150 316350
rect 565218 316294 565274 316350
rect 565342 316294 565398 316350
rect 564970 316170 565026 316226
rect 565094 316170 565150 316226
rect 565218 316170 565274 316226
rect 565342 316170 565398 316226
rect 564970 316046 565026 316102
rect 565094 316046 565150 316102
rect 565218 316046 565274 316102
rect 565342 316046 565398 316102
rect 564970 315922 565026 315978
rect 565094 315922 565150 315978
rect 565218 315922 565274 315978
rect 565342 315922 565398 315978
rect 564970 298294 565026 298350
rect 565094 298294 565150 298350
rect 565218 298294 565274 298350
rect 565342 298294 565398 298350
rect 564970 298170 565026 298226
rect 565094 298170 565150 298226
rect 565218 298170 565274 298226
rect 565342 298170 565398 298226
rect 564970 298046 565026 298102
rect 565094 298046 565150 298102
rect 565218 298046 565274 298102
rect 565342 298046 565398 298102
rect 564970 297922 565026 297978
rect 565094 297922 565150 297978
rect 565218 297922 565274 297978
rect 565342 297922 565398 297978
rect 564970 280294 565026 280350
rect 565094 280294 565150 280350
rect 565218 280294 565274 280350
rect 565342 280294 565398 280350
rect 564970 280170 565026 280226
rect 565094 280170 565150 280226
rect 565218 280170 565274 280226
rect 565342 280170 565398 280226
rect 564970 280046 565026 280102
rect 565094 280046 565150 280102
rect 565218 280046 565274 280102
rect 565342 280046 565398 280102
rect 564970 279922 565026 279978
rect 565094 279922 565150 279978
rect 565218 279922 565274 279978
rect 565342 279922 565398 279978
rect 564970 262294 565026 262350
rect 565094 262294 565150 262350
rect 565218 262294 565274 262350
rect 565342 262294 565398 262350
rect 564970 262170 565026 262226
rect 565094 262170 565150 262226
rect 565218 262170 565274 262226
rect 565342 262170 565398 262226
rect 564970 262046 565026 262102
rect 565094 262046 565150 262102
rect 565218 262046 565274 262102
rect 565342 262046 565398 262102
rect 564970 261922 565026 261978
rect 565094 261922 565150 261978
rect 565218 261922 565274 261978
rect 565342 261922 565398 261978
rect 564970 244294 565026 244350
rect 565094 244294 565150 244350
rect 565218 244294 565274 244350
rect 565342 244294 565398 244350
rect 564970 244170 565026 244226
rect 565094 244170 565150 244226
rect 565218 244170 565274 244226
rect 565342 244170 565398 244226
rect 564970 244046 565026 244102
rect 565094 244046 565150 244102
rect 565218 244046 565274 244102
rect 565342 244046 565398 244102
rect 564970 243922 565026 243978
rect 565094 243922 565150 243978
rect 565218 243922 565274 243978
rect 565342 243922 565398 243978
rect 564970 226294 565026 226350
rect 565094 226294 565150 226350
rect 565218 226294 565274 226350
rect 565342 226294 565398 226350
rect 564970 226170 565026 226226
rect 565094 226170 565150 226226
rect 565218 226170 565274 226226
rect 565342 226170 565398 226226
rect 564970 226046 565026 226102
rect 565094 226046 565150 226102
rect 565218 226046 565274 226102
rect 565342 226046 565398 226102
rect 564970 225922 565026 225978
rect 565094 225922 565150 225978
rect 565218 225922 565274 225978
rect 565342 225922 565398 225978
rect 564970 208294 565026 208350
rect 565094 208294 565150 208350
rect 565218 208294 565274 208350
rect 565342 208294 565398 208350
rect 564970 208170 565026 208226
rect 565094 208170 565150 208226
rect 565218 208170 565274 208226
rect 565342 208170 565398 208226
rect 564970 208046 565026 208102
rect 565094 208046 565150 208102
rect 565218 208046 565274 208102
rect 565342 208046 565398 208102
rect 564970 207922 565026 207978
rect 565094 207922 565150 207978
rect 565218 207922 565274 207978
rect 565342 207922 565398 207978
rect 564970 190294 565026 190350
rect 565094 190294 565150 190350
rect 565218 190294 565274 190350
rect 565342 190294 565398 190350
rect 564970 190170 565026 190226
rect 565094 190170 565150 190226
rect 565218 190170 565274 190226
rect 565342 190170 565398 190226
rect 564970 190046 565026 190102
rect 565094 190046 565150 190102
rect 565218 190046 565274 190102
rect 565342 190046 565398 190102
rect 564970 189922 565026 189978
rect 565094 189922 565150 189978
rect 565218 189922 565274 189978
rect 565342 189922 565398 189978
rect 564970 172294 565026 172350
rect 565094 172294 565150 172350
rect 565218 172294 565274 172350
rect 565342 172294 565398 172350
rect 564970 172170 565026 172226
rect 565094 172170 565150 172226
rect 565218 172170 565274 172226
rect 565342 172170 565398 172226
rect 564970 172046 565026 172102
rect 565094 172046 565150 172102
rect 565218 172046 565274 172102
rect 565342 172046 565398 172102
rect 564970 171922 565026 171978
rect 565094 171922 565150 171978
rect 565218 171922 565274 171978
rect 565342 171922 565398 171978
rect 564970 154294 565026 154350
rect 565094 154294 565150 154350
rect 565218 154294 565274 154350
rect 565342 154294 565398 154350
rect 564970 154170 565026 154226
rect 565094 154170 565150 154226
rect 565218 154170 565274 154226
rect 565342 154170 565398 154226
rect 564970 154046 565026 154102
rect 565094 154046 565150 154102
rect 565218 154046 565274 154102
rect 565342 154046 565398 154102
rect 564970 153922 565026 153978
rect 565094 153922 565150 153978
rect 565218 153922 565274 153978
rect 565342 153922 565398 153978
rect 564970 136294 565026 136350
rect 565094 136294 565150 136350
rect 565218 136294 565274 136350
rect 565342 136294 565398 136350
rect 564970 136170 565026 136226
rect 565094 136170 565150 136226
rect 565218 136170 565274 136226
rect 565342 136170 565398 136226
rect 564970 136046 565026 136102
rect 565094 136046 565150 136102
rect 565218 136046 565274 136102
rect 565342 136046 565398 136102
rect 564970 135922 565026 135978
rect 565094 135922 565150 135978
rect 565218 135922 565274 135978
rect 565342 135922 565398 135978
rect 564970 118294 565026 118350
rect 565094 118294 565150 118350
rect 565218 118294 565274 118350
rect 565342 118294 565398 118350
rect 564970 118170 565026 118226
rect 565094 118170 565150 118226
rect 565218 118170 565274 118226
rect 565342 118170 565398 118226
rect 564970 118046 565026 118102
rect 565094 118046 565150 118102
rect 565218 118046 565274 118102
rect 565342 118046 565398 118102
rect 564970 117922 565026 117978
rect 565094 117922 565150 117978
rect 565218 117922 565274 117978
rect 565342 117922 565398 117978
rect 564970 100294 565026 100350
rect 565094 100294 565150 100350
rect 565218 100294 565274 100350
rect 565342 100294 565398 100350
rect 564970 100170 565026 100226
rect 565094 100170 565150 100226
rect 565218 100170 565274 100226
rect 565342 100170 565398 100226
rect 564970 100046 565026 100102
rect 565094 100046 565150 100102
rect 565218 100046 565274 100102
rect 565342 100046 565398 100102
rect 564970 99922 565026 99978
rect 565094 99922 565150 99978
rect 565218 99922 565274 99978
rect 565342 99922 565398 99978
rect 564970 82294 565026 82350
rect 565094 82294 565150 82350
rect 565218 82294 565274 82350
rect 565342 82294 565398 82350
rect 564970 82170 565026 82226
rect 565094 82170 565150 82226
rect 565218 82170 565274 82226
rect 565342 82170 565398 82226
rect 564970 82046 565026 82102
rect 565094 82046 565150 82102
rect 565218 82046 565274 82102
rect 565342 82046 565398 82102
rect 564970 81922 565026 81978
rect 565094 81922 565150 81978
rect 565218 81922 565274 81978
rect 565342 81922 565398 81978
rect 564970 64294 565026 64350
rect 565094 64294 565150 64350
rect 565218 64294 565274 64350
rect 565342 64294 565398 64350
rect 564970 64170 565026 64226
rect 565094 64170 565150 64226
rect 565218 64170 565274 64226
rect 565342 64170 565398 64226
rect 564970 64046 565026 64102
rect 565094 64046 565150 64102
rect 565218 64046 565274 64102
rect 565342 64046 565398 64102
rect 564970 63922 565026 63978
rect 565094 63922 565150 63978
rect 565218 63922 565274 63978
rect 565342 63922 565398 63978
rect 564970 46294 565026 46350
rect 565094 46294 565150 46350
rect 565218 46294 565274 46350
rect 565342 46294 565398 46350
rect 564970 46170 565026 46226
rect 565094 46170 565150 46226
rect 565218 46170 565274 46226
rect 565342 46170 565398 46226
rect 564970 46046 565026 46102
rect 565094 46046 565150 46102
rect 565218 46046 565274 46102
rect 565342 46046 565398 46102
rect 564970 45922 565026 45978
rect 565094 45922 565150 45978
rect 565218 45922 565274 45978
rect 565342 45922 565398 45978
rect 564970 28294 565026 28350
rect 565094 28294 565150 28350
rect 565218 28294 565274 28350
rect 565342 28294 565398 28350
rect 564970 28170 565026 28226
rect 565094 28170 565150 28226
rect 565218 28170 565274 28226
rect 565342 28170 565398 28226
rect 564970 28046 565026 28102
rect 565094 28046 565150 28102
rect 565218 28046 565274 28102
rect 565342 28046 565398 28102
rect 564970 27922 565026 27978
rect 565094 27922 565150 27978
rect 565218 27922 565274 27978
rect 565342 27922 565398 27978
rect 564970 10294 565026 10350
rect 565094 10294 565150 10350
rect 565218 10294 565274 10350
rect 565342 10294 565398 10350
rect 564970 10170 565026 10226
rect 565094 10170 565150 10226
rect 565218 10170 565274 10226
rect 565342 10170 565398 10226
rect 564970 10046 565026 10102
rect 565094 10046 565150 10102
rect 565218 10046 565274 10102
rect 565342 10046 565398 10102
rect 564970 9922 565026 9978
rect 565094 9922 565150 9978
rect 565218 9922 565274 9978
rect 565342 9922 565398 9978
rect 564970 -1176 565026 -1120
rect 565094 -1176 565150 -1120
rect 565218 -1176 565274 -1120
rect 565342 -1176 565398 -1120
rect 564970 -1300 565026 -1244
rect 565094 -1300 565150 -1244
rect 565218 -1300 565274 -1244
rect 565342 -1300 565398 -1244
rect 564970 -1424 565026 -1368
rect 565094 -1424 565150 -1368
rect 565218 -1424 565274 -1368
rect 565342 -1424 565398 -1368
rect 564970 -1548 565026 -1492
rect 565094 -1548 565150 -1492
rect 565218 -1548 565274 -1492
rect 565342 -1548 565398 -1492
rect 579250 597156 579306 597212
rect 579374 597156 579430 597212
rect 579498 597156 579554 597212
rect 579622 597156 579678 597212
rect 579250 597032 579306 597088
rect 579374 597032 579430 597088
rect 579498 597032 579554 597088
rect 579622 597032 579678 597088
rect 579250 596908 579306 596964
rect 579374 596908 579430 596964
rect 579498 596908 579554 596964
rect 579622 596908 579678 596964
rect 579250 596784 579306 596840
rect 579374 596784 579430 596840
rect 579498 596784 579554 596840
rect 579622 596784 579678 596840
rect 579250 580294 579306 580350
rect 579374 580294 579430 580350
rect 579498 580294 579554 580350
rect 579622 580294 579678 580350
rect 579250 580170 579306 580226
rect 579374 580170 579430 580226
rect 579498 580170 579554 580226
rect 579622 580170 579678 580226
rect 579250 580046 579306 580102
rect 579374 580046 579430 580102
rect 579498 580046 579554 580102
rect 579622 580046 579678 580102
rect 579250 579922 579306 579978
rect 579374 579922 579430 579978
rect 579498 579922 579554 579978
rect 579622 579922 579678 579978
rect 579250 562294 579306 562350
rect 579374 562294 579430 562350
rect 579498 562294 579554 562350
rect 579622 562294 579678 562350
rect 579250 562170 579306 562226
rect 579374 562170 579430 562226
rect 579498 562170 579554 562226
rect 579622 562170 579678 562226
rect 579250 562046 579306 562102
rect 579374 562046 579430 562102
rect 579498 562046 579554 562102
rect 579622 562046 579678 562102
rect 579250 561922 579306 561978
rect 579374 561922 579430 561978
rect 579498 561922 579554 561978
rect 579622 561922 579678 561978
rect 579250 544294 579306 544350
rect 579374 544294 579430 544350
rect 579498 544294 579554 544350
rect 579622 544294 579678 544350
rect 579250 544170 579306 544226
rect 579374 544170 579430 544226
rect 579498 544170 579554 544226
rect 579622 544170 579678 544226
rect 579250 544046 579306 544102
rect 579374 544046 579430 544102
rect 579498 544046 579554 544102
rect 579622 544046 579678 544102
rect 579250 543922 579306 543978
rect 579374 543922 579430 543978
rect 579498 543922 579554 543978
rect 579622 543922 579678 543978
rect 579250 526294 579306 526350
rect 579374 526294 579430 526350
rect 579498 526294 579554 526350
rect 579622 526294 579678 526350
rect 579250 526170 579306 526226
rect 579374 526170 579430 526226
rect 579498 526170 579554 526226
rect 579622 526170 579678 526226
rect 579250 526046 579306 526102
rect 579374 526046 579430 526102
rect 579498 526046 579554 526102
rect 579622 526046 579678 526102
rect 579250 525922 579306 525978
rect 579374 525922 579430 525978
rect 579498 525922 579554 525978
rect 579622 525922 579678 525978
rect 579250 508294 579306 508350
rect 579374 508294 579430 508350
rect 579498 508294 579554 508350
rect 579622 508294 579678 508350
rect 579250 508170 579306 508226
rect 579374 508170 579430 508226
rect 579498 508170 579554 508226
rect 579622 508170 579678 508226
rect 579250 508046 579306 508102
rect 579374 508046 579430 508102
rect 579498 508046 579554 508102
rect 579622 508046 579678 508102
rect 579250 507922 579306 507978
rect 579374 507922 579430 507978
rect 579498 507922 579554 507978
rect 579622 507922 579678 507978
rect 579250 490294 579306 490350
rect 579374 490294 579430 490350
rect 579498 490294 579554 490350
rect 579622 490294 579678 490350
rect 579250 490170 579306 490226
rect 579374 490170 579430 490226
rect 579498 490170 579554 490226
rect 579622 490170 579678 490226
rect 579250 490046 579306 490102
rect 579374 490046 579430 490102
rect 579498 490046 579554 490102
rect 579622 490046 579678 490102
rect 579250 489922 579306 489978
rect 579374 489922 579430 489978
rect 579498 489922 579554 489978
rect 579622 489922 579678 489978
rect 579250 472294 579306 472350
rect 579374 472294 579430 472350
rect 579498 472294 579554 472350
rect 579622 472294 579678 472350
rect 579250 472170 579306 472226
rect 579374 472170 579430 472226
rect 579498 472170 579554 472226
rect 579622 472170 579678 472226
rect 579250 472046 579306 472102
rect 579374 472046 579430 472102
rect 579498 472046 579554 472102
rect 579622 472046 579678 472102
rect 579250 471922 579306 471978
rect 579374 471922 579430 471978
rect 579498 471922 579554 471978
rect 579622 471922 579678 471978
rect 579250 454294 579306 454350
rect 579374 454294 579430 454350
rect 579498 454294 579554 454350
rect 579622 454294 579678 454350
rect 579250 454170 579306 454226
rect 579374 454170 579430 454226
rect 579498 454170 579554 454226
rect 579622 454170 579678 454226
rect 579250 454046 579306 454102
rect 579374 454046 579430 454102
rect 579498 454046 579554 454102
rect 579622 454046 579678 454102
rect 579250 453922 579306 453978
rect 579374 453922 579430 453978
rect 579498 453922 579554 453978
rect 579622 453922 579678 453978
rect 579250 436294 579306 436350
rect 579374 436294 579430 436350
rect 579498 436294 579554 436350
rect 579622 436294 579678 436350
rect 579250 436170 579306 436226
rect 579374 436170 579430 436226
rect 579498 436170 579554 436226
rect 579622 436170 579678 436226
rect 579250 436046 579306 436102
rect 579374 436046 579430 436102
rect 579498 436046 579554 436102
rect 579622 436046 579678 436102
rect 579250 435922 579306 435978
rect 579374 435922 579430 435978
rect 579498 435922 579554 435978
rect 579622 435922 579678 435978
rect 579250 418294 579306 418350
rect 579374 418294 579430 418350
rect 579498 418294 579554 418350
rect 579622 418294 579678 418350
rect 579250 418170 579306 418226
rect 579374 418170 579430 418226
rect 579498 418170 579554 418226
rect 579622 418170 579678 418226
rect 579250 418046 579306 418102
rect 579374 418046 579430 418102
rect 579498 418046 579554 418102
rect 579622 418046 579678 418102
rect 579250 417922 579306 417978
rect 579374 417922 579430 417978
rect 579498 417922 579554 417978
rect 579622 417922 579678 417978
rect 579250 400294 579306 400350
rect 579374 400294 579430 400350
rect 579498 400294 579554 400350
rect 579622 400294 579678 400350
rect 579250 400170 579306 400226
rect 579374 400170 579430 400226
rect 579498 400170 579554 400226
rect 579622 400170 579678 400226
rect 579250 400046 579306 400102
rect 579374 400046 579430 400102
rect 579498 400046 579554 400102
rect 579622 400046 579678 400102
rect 579250 399922 579306 399978
rect 579374 399922 579430 399978
rect 579498 399922 579554 399978
rect 579622 399922 579678 399978
rect 579250 382294 579306 382350
rect 579374 382294 579430 382350
rect 579498 382294 579554 382350
rect 579622 382294 579678 382350
rect 579250 382170 579306 382226
rect 579374 382170 579430 382226
rect 579498 382170 579554 382226
rect 579622 382170 579678 382226
rect 579250 382046 579306 382102
rect 579374 382046 579430 382102
rect 579498 382046 579554 382102
rect 579622 382046 579678 382102
rect 579250 381922 579306 381978
rect 579374 381922 579430 381978
rect 579498 381922 579554 381978
rect 579622 381922 579678 381978
rect 579250 364294 579306 364350
rect 579374 364294 579430 364350
rect 579498 364294 579554 364350
rect 579622 364294 579678 364350
rect 579250 364170 579306 364226
rect 579374 364170 579430 364226
rect 579498 364170 579554 364226
rect 579622 364170 579678 364226
rect 579250 364046 579306 364102
rect 579374 364046 579430 364102
rect 579498 364046 579554 364102
rect 579622 364046 579678 364102
rect 579250 363922 579306 363978
rect 579374 363922 579430 363978
rect 579498 363922 579554 363978
rect 579622 363922 579678 363978
rect 579250 346294 579306 346350
rect 579374 346294 579430 346350
rect 579498 346294 579554 346350
rect 579622 346294 579678 346350
rect 579250 346170 579306 346226
rect 579374 346170 579430 346226
rect 579498 346170 579554 346226
rect 579622 346170 579678 346226
rect 579250 346046 579306 346102
rect 579374 346046 579430 346102
rect 579498 346046 579554 346102
rect 579622 346046 579678 346102
rect 579250 345922 579306 345978
rect 579374 345922 579430 345978
rect 579498 345922 579554 345978
rect 579622 345922 579678 345978
rect 579250 328294 579306 328350
rect 579374 328294 579430 328350
rect 579498 328294 579554 328350
rect 579622 328294 579678 328350
rect 579250 328170 579306 328226
rect 579374 328170 579430 328226
rect 579498 328170 579554 328226
rect 579622 328170 579678 328226
rect 579250 328046 579306 328102
rect 579374 328046 579430 328102
rect 579498 328046 579554 328102
rect 579622 328046 579678 328102
rect 579250 327922 579306 327978
rect 579374 327922 579430 327978
rect 579498 327922 579554 327978
rect 579622 327922 579678 327978
rect 579250 310294 579306 310350
rect 579374 310294 579430 310350
rect 579498 310294 579554 310350
rect 579622 310294 579678 310350
rect 579250 310170 579306 310226
rect 579374 310170 579430 310226
rect 579498 310170 579554 310226
rect 579622 310170 579678 310226
rect 579250 310046 579306 310102
rect 579374 310046 579430 310102
rect 579498 310046 579554 310102
rect 579622 310046 579678 310102
rect 579250 309922 579306 309978
rect 579374 309922 579430 309978
rect 579498 309922 579554 309978
rect 579622 309922 579678 309978
rect 579250 292294 579306 292350
rect 579374 292294 579430 292350
rect 579498 292294 579554 292350
rect 579622 292294 579678 292350
rect 579250 292170 579306 292226
rect 579374 292170 579430 292226
rect 579498 292170 579554 292226
rect 579622 292170 579678 292226
rect 579250 292046 579306 292102
rect 579374 292046 579430 292102
rect 579498 292046 579554 292102
rect 579622 292046 579678 292102
rect 579250 291922 579306 291978
rect 579374 291922 579430 291978
rect 579498 291922 579554 291978
rect 579622 291922 579678 291978
rect 579250 274294 579306 274350
rect 579374 274294 579430 274350
rect 579498 274294 579554 274350
rect 579622 274294 579678 274350
rect 579250 274170 579306 274226
rect 579374 274170 579430 274226
rect 579498 274170 579554 274226
rect 579622 274170 579678 274226
rect 579250 274046 579306 274102
rect 579374 274046 579430 274102
rect 579498 274046 579554 274102
rect 579622 274046 579678 274102
rect 579250 273922 579306 273978
rect 579374 273922 579430 273978
rect 579498 273922 579554 273978
rect 579622 273922 579678 273978
rect 579250 256294 579306 256350
rect 579374 256294 579430 256350
rect 579498 256294 579554 256350
rect 579622 256294 579678 256350
rect 579250 256170 579306 256226
rect 579374 256170 579430 256226
rect 579498 256170 579554 256226
rect 579622 256170 579678 256226
rect 579250 256046 579306 256102
rect 579374 256046 579430 256102
rect 579498 256046 579554 256102
rect 579622 256046 579678 256102
rect 579250 255922 579306 255978
rect 579374 255922 579430 255978
rect 579498 255922 579554 255978
rect 579622 255922 579678 255978
rect 579250 238294 579306 238350
rect 579374 238294 579430 238350
rect 579498 238294 579554 238350
rect 579622 238294 579678 238350
rect 579250 238170 579306 238226
rect 579374 238170 579430 238226
rect 579498 238170 579554 238226
rect 579622 238170 579678 238226
rect 579250 238046 579306 238102
rect 579374 238046 579430 238102
rect 579498 238046 579554 238102
rect 579622 238046 579678 238102
rect 579250 237922 579306 237978
rect 579374 237922 579430 237978
rect 579498 237922 579554 237978
rect 579622 237922 579678 237978
rect 579250 220294 579306 220350
rect 579374 220294 579430 220350
rect 579498 220294 579554 220350
rect 579622 220294 579678 220350
rect 579250 220170 579306 220226
rect 579374 220170 579430 220226
rect 579498 220170 579554 220226
rect 579622 220170 579678 220226
rect 579250 220046 579306 220102
rect 579374 220046 579430 220102
rect 579498 220046 579554 220102
rect 579622 220046 579678 220102
rect 579250 219922 579306 219978
rect 579374 219922 579430 219978
rect 579498 219922 579554 219978
rect 579622 219922 579678 219978
rect 579250 202294 579306 202350
rect 579374 202294 579430 202350
rect 579498 202294 579554 202350
rect 579622 202294 579678 202350
rect 579250 202170 579306 202226
rect 579374 202170 579430 202226
rect 579498 202170 579554 202226
rect 579622 202170 579678 202226
rect 579250 202046 579306 202102
rect 579374 202046 579430 202102
rect 579498 202046 579554 202102
rect 579622 202046 579678 202102
rect 579250 201922 579306 201978
rect 579374 201922 579430 201978
rect 579498 201922 579554 201978
rect 579622 201922 579678 201978
rect 579250 184294 579306 184350
rect 579374 184294 579430 184350
rect 579498 184294 579554 184350
rect 579622 184294 579678 184350
rect 579250 184170 579306 184226
rect 579374 184170 579430 184226
rect 579498 184170 579554 184226
rect 579622 184170 579678 184226
rect 579250 184046 579306 184102
rect 579374 184046 579430 184102
rect 579498 184046 579554 184102
rect 579622 184046 579678 184102
rect 579250 183922 579306 183978
rect 579374 183922 579430 183978
rect 579498 183922 579554 183978
rect 579622 183922 579678 183978
rect 579250 166294 579306 166350
rect 579374 166294 579430 166350
rect 579498 166294 579554 166350
rect 579622 166294 579678 166350
rect 579250 166170 579306 166226
rect 579374 166170 579430 166226
rect 579498 166170 579554 166226
rect 579622 166170 579678 166226
rect 579250 166046 579306 166102
rect 579374 166046 579430 166102
rect 579498 166046 579554 166102
rect 579622 166046 579678 166102
rect 579250 165922 579306 165978
rect 579374 165922 579430 165978
rect 579498 165922 579554 165978
rect 579622 165922 579678 165978
rect 579250 148294 579306 148350
rect 579374 148294 579430 148350
rect 579498 148294 579554 148350
rect 579622 148294 579678 148350
rect 579250 148170 579306 148226
rect 579374 148170 579430 148226
rect 579498 148170 579554 148226
rect 579622 148170 579678 148226
rect 579250 148046 579306 148102
rect 579374 148046 579430 148102
rect 579498 148046 579554 148102
rect 579622 148046 579678 148102
rect 579250 147922 579306 147978
rect 579374 147922 579430 147978
rect 579498 147922 579554 147978
rect 579622 147922 579678 147978
rect 579250 130294 579306 130350
rect 579374 130294 579430 130350
rect 579498 130294 579554 130350
rect 579622 130294 579678 130350
rect 579250 130170 579306 130226
rect 579374 130170 579430 130226
rect 579498 130170 579554 130226
rect 579622 130170 579678 130226
rect 579250 130046 579306 130102
rect 579374 130046 579430 130102
rect 579498 130046 579554 130102
rect 579622 130046 579678 130102
rect 579250 129922 579306 129978
rect 579374 129922 579430 129978
rect 579498 129922 579554 129978
rect 579622 129922 579678 129978
rect 579250 112294 579306 112350
rect 579374 112294 579430 112350
rect 579498 112294 579554 112350
rect 579622 112294 579678 112350
rect 579250 112170 579306 112226
rect 579374 112170 579430 112226
rect 579498 112170 579554 112226
rect 579622 112170 579678 112226
rect 579250 112046 579306 112102
rect 579374 112046 579430 112102
rect 579498 112046 579554 112102
rect 579622 112046 579678 112102
rect 579250 111922 579306 111978
rect 579374 111922 579430 111978
rect 579498 111922 579554 111978
rect 579622 111922 579678 111978
rect 579250 94294 579306 94350
rect 579374 94294 579430 94350
rect 579498 94294 579554 94350
rect 579622 94294 579678 94350
rect 579250 94170 579306 94226
rect 579374 94170 579430 94226
rect 579498 94170 579554 94226
rect 579622 94170 579678 94226
rect 579250 94046 579306 94102
rect 579374 94046 579430 94102
rect 579498 94046 579554 94102
rect 579622 94046 579678 94102
rect 579250 93922 579306 93978
rect 579374 93922 579430 93978
rect 579498 93922 579554 93978
rect 579622 93922 579678 93978
rect 579250 76294 579306 76350
rect 579374 76294 579430 76350
rect 579498 76294 579554 76350
rect 579622 76294 579678 76350
rect 579250 76170 579306 76226
rect 579374 76170 579430 76226
rect 579498 76170 579554 76226
rect 579622 76170 579678 76226
rect 579250 76046 579306 76102
rect 579374 76046 579430 76102
rect 579498 76046 579554 76102
rect 579622 76046 579678 76102
rect 579250 75922 579306 75978
rect 579374 75922 579430 75978
rect 579498 75922 579554 75978
rect 579622 75922 579678 75978
rect 579250 58294 579306 58350
rect 579374 58294 579430 58350
rect 579498 58294 579554 58350
rect 579622 58294 579678 58350
rect 579250 58170 579306 58226
rect 579374 58170 579430 58226
rect 579498 58170 579554 58226
rect 579622 58170 579678 58226
rect 579250 58046 579306 58102
rect 579374 58046 579430 58102
rect 579498 58046 579554 58102
rect 579622 58046 579678 58102
rect 579250 57922 579306 57978
rect 579374 57922 579430 57978
rect 579498 57922 579554 57978
rect 579622 57922 579678 57978
rect 579250 40294 579306 40350
rect 579374 40294 579430 40350
rect 579498 40294 579554 40350
rect 579622 40294 579678 40350
rect 579250 40170 579306 40226
rect 579374 40170 579430 40226
rect 579498 40170 579554 40226
rect 579622 40170 579678 40226
rect 579250 40046 579306 40102
rect 579374 40046 579430 40102
rect 579498 40046 579554 40102
rect 579622 40046 579678 40102
rect 579250 39922 579306 39978
rect 579374 39922 579430 39978
rect 579498 39922 579554 39978
rect 579622 39922 579678 39978
rect 579250 22294 579306 22350
rect 579374 22294 579430 22350
rect 579498 22294 579554 22350
rect 579622 22294 579678 22350
rect 579250 22170 579306 22226
rect 579374 22170 579430 22226
rect 579498 22170 579554 22226
rect 579622 22170 579678 22226
rect 579250 22046 579306 22102
rect 579374 22046 579430 22102
rect 579498 22046 579554 22102
rect 579622 22046 579678 22102
rect 579250 21922 579306 21978
rect 579374 21922 579430 21978
rect 579498 21922 579554 21978
rect 579622 21922 579678 21978
rect 579250 4294 579306 4350
rect 579374 4294 579430 4350
rect 579498 4294 579554 4350
rect 579622 4294 579678 4350
rect 579250 4170 579306 4226
rect 579374 4170 579430 4226
rect 579498 4170 579554 4226
rect 579622 4170 579678 4226
rect 579250 4046 579306 4102
rect 579374 4046 579430 4102
rect 579498 4046 579554 4102
rect 579622 4046 579678 4102
rect 579250 3922 579306 3978
rect 579374 3922 579430 3978
rect 579498 3922 579554 3978
rect 579622 3922 579678 3978
rect 579250 -216 579306 -160
rect 579374 -216 579430 -160
rect 579498 -216 579554 -160
rect 579622 -216 579678 -160
rect 579250 -340 579306 -284
rect 579374 -340 579430 -284
rect 579498 -340 579554 -284
rect 579622 -340 579678 -284
rect 579250 -464 579306 -408
rect 579374 -464 579430 -408
rect 579498 -464 579554 -408
rect 579622 -464 579678 -408
rect 579250 -588 579306 -532
rect 579374 -588 579430 -532
rect 579498 -588 579554 -532
rect 579622 -588 579678 -532
rect 582970 598116 583026 598172
rect 583094 598116 583150 598172
rect 583218 598116 583274 598172
rect 583342 598116 583398 598172
rect 582970 597992 583026 598048
rect 583094 597992 583150 598048
rect 583218 597992 583274 598048
rect 583342 597992 583398 598048
rect 582970 597868 583026 597924
rect 583094 597868 583150 597924
rect 583218 597868 583274 597924
rect 583342 597868 583398 597924
rect 582970 597744 583026 597800
rect 583094 597744 583150 597800
rect 583218 597744 583274 597800
rect 583342 597744 583398 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 582970 586294 583026 586350
rect 583094 586294 583150 586350
rect 583218 586294 583274 586350
rect 583342 586294 583398 586350
rect 582970 586170 583026 586226
rect 583094 586170 583150 586226
rect 583218 586170 583274 586226
rect 583342 586170 583398 586226
rect 582970 586046 583026 586102
rect 583094 586046 583150 586102
rect 583218 586046 583274 586102
rect 583342 586046 583398 586102
rect 582970 585922 583026 585978
rect 583094 585922 583150 585978
rect 583218 585922 583274 585978
rect 583342 585922 583398 585978
rect 582970 568294 583026 568350
rect 583094 568294 583150 568350
rect 583218 568294 583274 568350
rect 583342 568294 583398 568350
rect 582970 568170 583026 568226
rect 583094 568170 583150 568226
rect 583218 568170 583274 568226
rect 583342 568170 583398 568226
rect 582970 568046 583026 568102
rect 583094 568046 583150 568102
rect 583218 568046 583274 568102
rect 583342 568046 583398 568102
rect 582970 567922 583026 567978
rect 583094 567922 583150 567978
rect 583218 567922 583274 567978
rect 583342 567922 583398 567978
rect 582970 550294 583026 550350
rect 583094 550294 583150 550350
rect 583218 550294 583274 550350
rect 583342 550294 583398 550350
rect 582970 550170 583026 550226
rect 583094 550170 583150 550226
rect 583218 550170 583274 550226
rect 583342 550170 583398 550226
rect 582970 550046 583026 550102
rect 583094 550046 583150 550102
rect 583218 550046 583274 550102
rect 583342 550046 583398 550102
rect 582970 549922 583026 549978
rect 583094 549922 583150 549978
rect 583218 549922 583274 549978
rect 583342 549922 583398 549978
rect 582970 532294 583026 532350
rect 583094 532294 583150 532350
rect 583218 532294 583274 532350
rect 583342 532294 583398 532350
rect 582970 532170 583026 532226
rect 583094 532170 583150 532226
rect 583218 532170 583274 532226
rect 583342 532170 583398 532226
rect 582970 532046 583026 532102
rect 583094 532046 583150 532102
rect 583218 532046 583274 532102
rect 583342 532046 583398 532102
rect 582970 531922 583026 531978
rect 583094 531922 583150 531978
rect 583218 531922 583274 531978
rect 583342 531922 583398 531978
rect 582970 514294 583026 514350
rect 583094 514294 583150 514350
rect 583218 514294 583274 514350
rect 583342 514294 583398 514350
rect 582970 514170 583026 514226
rect 583094 514170 583150 514226
rect 583218 514170 583274 514226
rect 583342 514170 583398 514226
rect 582970 514046 583026 514102
rect 583094 514046 583150 514102
rect 583218 514046 583274 514102
rect 583342 514046 583398 514102
rect 582970 513922 583026 513978
rect 583094 513922 583150 513978
rect 583218 513922 583274 513978
rect 583342 513922 583398 513978
rect 582970 496294 583026 496350
rect 583094 496294 583150 496350
rect 583218 496294 583274 496350
rect 583342 496294 583398 496350
rect 582970 496170 583026 496226
rect 583094 496170 583150 496226
rect 583218 496170 583274 496226
rect 583342 496170 583398 496226
rect 582970 496046 583026 496102
rect 583094 496046 583150 496102
rect 583218 496046 583274 496102
rect 583342 496046 583398 496102
rect 582970 495922 583026 495978
rect 583094 495922 583150 495978
rect 583218 495922 583274 495978
rect 583342 495922 583398 495978
rect 582970 478294 583026 478350
rect 583094 478294 583150 478350
rect 583218 478294 583274 478350
rect 583342 478294 583398 478350
rect 582970 478170 583026 478226
rect 583094 478170 583150 478226
rect 583218 478170 583274 478226
rect 583342 478170 583398 478226
rect 582970 478046 583026 478102
rect 583094 478046 583150 478102
rect 583218 478046 583274 478102
rect 583342 478046 583398 478102
rect 582970 477922 583026 477978
rect 583094 477922 583150 477978
rect 583218 477922 583274 477978
rect 583342 477922 583398 477978
rect 582970 460294 583026 460350
rect 583094 460294 583150 460350
rect 583218 460294 583274 460350
rect 583342 460294 583398 460350
rect 582970 460170 583026 460226
rect 583094 460170 583150 460226
rect 583218 460170 583274 460226
rect 583342 460170 583398 460226
rect 582970 460046 583026 460102
rect 583094 460046 583150 460102
rect 583218 460046 583274 460102
rect 583342 460046 583398 460102
rect 582970 459922 583026 459978
rect 583094 459922 583150 459978
rect 583218 459922 583274 459978
rect 583342 459922 583398 459978
rect 582970 442294 583026 442350
rect 583094 442294 583150 442350
rect 583218 442294 583274 442350
rect 583342 442294 583398 442350
rect 582970 442170 583026 442226
rect 583094 442170 583150 442226
rect 583218 442170 583274 442226
rect 583342 442170 583398 442226
rect 582970 442046 583026 442102
rect 583094 442046 583150 442102
rect 583218 442046 583274 442102
rect 583342 442046 583398 442102
rect 582970 441922 583026 441978
rect 583094 441922 583150 441978
rect 583218 441922 583274 441978
rect 583342 441922 583398 441978
rect 582970 424294 583026 424350
rect 583094 424294 583150 424350
rect 583218 424294 583274 424350
rect 583342 424294 583398 424350
rect 582970 424170 583026 424226
rect 583094 424170 583150 424226
rect 583218 424170 583274 424226
rect 583342 424170 583398 424226
rect 582970 424046 583026 424102
rect 583094 424046 583150 424102
rect 583218 424046 583274 424102
rect 583342 424046 583398 424102
rect 582970 423922 583026 423978
rect 583094 423922 583150 423978
rect 583218 423922 583274 423978
rect 583342 423922 583398 423978
rect 582970 406294 583026 406350
rect 583094 406294 583150 406350
rect 583218 406294 583274 406350
rect 583342 406294 583398 406350
rect 582970 406170 583026 406226
rect 583094 406170 583150 406226
rect 583218 406170 583274 406226
rect 583342 406170 583398 406226
rect 582970 406046 583026 406102
rect 583094 406046 583150 406102
rect 583218 406046 583274 406102
rect 583342 406046 583398 406102
rect 582970 405922 583026 405978
rect 583094 405922 583150 405978
rect 583218 405922 583274 405978
rect 583342 405922 583398 405978
rect 582970 388294 583026 388350
rect 583094 388294 583150 388350
rect 583218 388294 583274 388350
rect 583342 388294 583398 388350
rect 582970 388170 583026 388226
rect 583094 388170 583150 388226
rect 583218 388170 583274 388226
rect 583342 388170 583398 388226
rect 582970 388046 583026 388102
rect 583094 388046 583150 388102
rect 583218 388046 583274 388102
rect 583342 388046 583398 388102
rect 582970 387922 583026 387978
rect 583094 387922 583150 387978
rect 583218 387922 583274 387978
rect 583342 387922 583398 387978
rect 582970 370294 583026 370350
rect 583094 370294 583150 370350
rect 583218 370294 583274 370350
rect 583342 370294 583398 370350
rect 582970 370170 583026 370226
rect 583094 370170 583150 370226
rect 583218 370170 583274 370226
rect 583342 370170 583398 370226
rect 582970 370046 583026 370102
rect 583094 370046 583150 370102
rect 583218 370046 583274 370102
rect 583342 370046 583398 370102
rect 582970 369922 583026 369978
rect 583094 369922 583150 369978
rect 583218 369922 583274 369978
rect 583342 369922 583398 369978
rect 582970 352294 583026 352350
rect 583094 352294 583150 352350
rect 583218 352294 583274 352350
rect 583342 352294 583398 352350
rect 582970 352170 583026 352226
rect 583094 352170 583150 352226
rect 583218 352170 583274 352226
rect 583342 352170 583398 352226
rect 582970 352046 583026 352102
rect 583094 352046 583150 352102
rect 583218 352046 583274 352102
rect 583342 352046 583398 352102
rect 582970 351922 583026 351978
rect 583094 351922 583150 351978
rect 583218 351922 583274 351978
rect 583342 351922 583398 351978
rect 582970 334294 583026 334350
rect 583094 334294 583150 334350
rect 583218 334294 583274 334350
rect 583342 334294 583398 334350
rect 582970 334170 583026 334226
rect 583094 334170 583150 334226
rect 583218 334170 583274 334226
rect 583342 334170 583398 334226
rect 582970 334046 583026 334102
rect 583094 334046 583150 334102
rect 583218 334046 583274 334102
rect 583342 334046 583398 334102
rect 582970 333922 583026 333978
rect 583094 333922 583150 333978
rect 583218 333922 583274 333978
rect 583342 333922 583398 333978
rect 582970 316294 583026 316350
rect 583094 316294 583150 316350
rect 583218 316294 583274 316350
rect 583342 316294 583398 316350
rect 582970 316170 583026 316226
rect 583094 316170 583150 316226
rect 583218 316170 583274 316226
rect 583342 316170 583398 316226
rect 582970 316046 583026 316102
rect 583094 316046 583150 316102
rect 583218 316046 583274 316102
rect 583342 316046 583398 316102
rect 582970 315922 583026 315978
rect 583094 315922 583150 315978
rect 583218 315922 583274 315978
rect 583342 315922 583398 315978
rect 582970 298294 583026 298350
rect 583094 298294 583150 298350
rect 583218 298294 583274 298350
rect 583342 298294 583398 298350
rect 582970 298170 583026 298226
rect 583094 298170 583150 298226
rect 583218 298170 583274 298226
rect 583342 298170 583398 298226
rect 582970 298046 583026 298102
rect 583094 298046 583150 298102
rect 583218 298046 583274 298102
rect 583342 298046 583398 298102
rect 582970 297922 583026 297978
rect 583094 297922 583150 297978
rect 583218 297922 583274 297978
rect 583342 297922 583398 297978
rect 582970 280294 583026 280350
rect 583094 280294 583150 280350
rect 583218 280294 583274 280350
rect 583342 280294 583398 280350
rect 582970 280170 583026 280226
rect 583094 280170 583150 280226
rect 583218 280170 583274 280226
rect 583342 280170 583398 280226
rect 582970 280046 583026 280102
rect 583094 280046 583150 280102
rect 583218 280046 583274 280102
rect 583342 280046 583398 280102
rect 582970 279922 583026 279978
rect 583094 279922 583150 279978
rect 583218 279922 583274 279978
rect 583342 279922 583398 279978
rect 582970 262294 583026 262350
rect 583094 262294 583150 262350
rect 583218 262294 583274 262350
rect 583342 262294 583398 262350
rect 582970 262170 583026 262226
rect 583094 262170 583150 262226
rect 583218 262170 583274 262226
rect 583342 262170 583398 262226
rect 582970 262046 583026 262102
rect 583094 262046 583150 262102
rect 583218 262046 583274 262102
rect 583342 262046 583398 262102
rect 582970 261922 583026 261978
rect 583094 261922 583150 261978
rect 583218 261922 583274 261978
rect 583342 261922 583398 261978
rect 582970 244294 583026 244350
rect 583094 244294 583150 244350
rect 583218 244294 583274 244350
rect 583342 244294 583398 244350
rect 582970 244170 583026 244226
rect 583094 244170 583150 244226
rect 583218 244170 583274 244226
rect 583342 244170 583398 244226
rect 582970 244046 583026 244102
rect 583094 244046 583150 244102
rect 583218 244046 583274 244102
rect 583342 244046 583398 244102
rect 582970 243922 583026 243978
rect 583094 243922 583150 243978
rect 583218 243922 583274 243978
rect 583342 243922 583398 243978
rect 582970 226294 583026 226350
rect 583094 226294 583150 226350
rect 583218 226294 583274 226350
rect 583342 226294 583398 226350
rect 582970 226170 583026 226226
rect 583094 226170 583150 226226
rect 583218 226170 583274 226226
rect 583342 226170 583398 226226
rect 582970 226046 583026 226102
rect 583094 226046 583150 226102
rect 583218 226046 583274 226102
rect 583342 226046 583398 226102
rect 582970 225922 583026 225978
rect 583094 225922 583150 225978
rect 583218 225922 583274 225978
rect 583342 225922 583398 225978
rect 582970 208294 583026 208350
rect 583094 208294 583150 208350
rect 583218 208294 583274 208350
rect 583342 208294 583398 208350
rect 582970 208170 583026 208226
rect 583094 208170 583150 208226
rect 583218 208170 583274 208226
rect 583342 208170 583398 208226
rect 582970 208046 583026 208102
rect 583094 208046 583150 208102
rect 583218 208046 583274 208102
rect 583342 208046 583398 208102
rect 582970 207922 583026 207978
rect 583094 207922 583150 207978
rect 583218 207922 583274 207978
rect 583342 207922 583398 207978
rect 582970 190294 583026 190350
rect 583094 190294 583150 190350
rect 583218 190294 583274 190350
rect 583342 190294 583398 190350
rect 582970 190170 583026 190226
rect 583094 190170 583150 190226
rect 583218 190170 583274 190226
rect 583342 190170 583398 190226
rect 582970 190046 583026 190102
rect 583094 190046 583150 190102
rect 583218 190046 583274 190102
rect 583342 190046 583398 190102
rect 582970 189922 583026 189978
rect 583094 189922 583150 189978
rect 583218 189922 583274 189978
rect 583342 189922 583398 189978
rect 582970 172294 583026 172350
rect 583094 172294 583150 172350
rect 583218 172294 583274 172350
rect 583342 172294 583398 172350
rect 582970 172170 583026 172226
rect 583094 172170 583150 172226
rect 583218 172170 583274 172226
rect 583342 172170 583398 172226
rect 582970 172046 583026 172102
rect 583094 172046 583150 172102
rect 583218 172046 583274 172102
rect 583342 172046 583398 172102
rect 582970 171922 583026 171978
rect 583094 171922 583150 171978
rect 583218 171922 583274 171978
rect 583342 171922 583398 171978
rect 582970 154294 583026 154350
rect 583094 154294 583150 154350
rect 583218 154294 583274 154350
rect 583342 154294 583398 154350
rect 582970 154170 583026 154226
rect 583094 154170 583150 154226
rect 583218 154170 583274 154226
rect 583342 154170 583398 154226
rect 582970 154046 583026 154102
rect 583094 154046 583150 154102
rect 583218 154046 583274 154102
rect 583342 154046 583398 154102
rect 582970 153922 583026 153978
rect 583094 153922 583150 153978
rect 583218 153922 583274 153978
rect 583342 153922 583398 153978
rect 582970 136294 583026 136350
rect 583094 136294 583150 136350
rect 583218 136294 583274 136350
rect 583342 136294 583398 136350
rect 582970 136170 583026 136226
rect 583094 136170 583150 136226
rect 583218 136170 583274 136226
rect 583342 136170 583398 136226
rect 582970 136046 583026 136102
rect 583094 136046 583150 136102
rect 583218 136046 583274 136102
rect 583342 136046 583398 136102
rect 582970 135922 583026 135978
rect 583094 135922 583150 135978
rect 583218 135922 583274 135978
rect 583342 135922 583398 135978
rect 582970 118294 583026 118350
rect 583094 118294 583150 118350
rect 583218 118294 583274 118350
rect 583342 118294 583398 118350
rect 582970 118170 583026 118226
rect 583094 118170 583150 118226
rect 583218 118170 583274 118226
rect 583342 118170 583398 118226
rect 582970 118046 583026 118102
rect 583094 118046 583150 118102
rect 583218 118046 583274 118102
rect 583342 118046 583398 118102
rect 582970 117922 583026 117978
rect 583094 117922 583150 117978
rect 583218 117922 583274 117978
rect 583342 117922 583398 117978
rect 582970 100294 583026 100350
rect 583094 100294 583150 100350
rect 583218 100294 583274 100350
rect 583342 100294 583398 100350
rect 582970 100170 583026 100226
rect 583094 100170 583150 100226
rect 583218 100170 583274 100226
rect 583342 100170 583398 100226
rect 582970 100046 583026 100102
rect 583094 100046 583150 100102
rect 583218 100046 583274 100102
rect 583342 100046 583398 100102
rect 582970 99922 583026 99978
rect 583094 99922 583150 99978
rect 583218 99922 583274 99978
rect 583342 99922 583398 99978
rect 582970 82294 583026 82350
rect 583094 82294 583150 82350
rect 583218 82294 583274 82350
rect 583342 82294 583398 82350
rect 582970 82170 583026 82226
rect 583094 82170 583150 82226
rect 583218 82170 583274 82226
rect 583342 82170 583398 82226
rect 582970 82046 583026 82102
rect 583094 82046 583150 82102
rect 583218 82046 583274 82102
rect 583342 82046 583398 82102
rect 582970 81922 583026 81978
rect 583094 81922 583150 81978
rect 583218 81922 583274 81978
rect 583342 81922 583398 81978
rect 582970 64294 583026 64350
rect 583094 64294 583150 64350
rect 583218 64294 583274 64350
rect 583342 64294 583398 64350
rect 582970 64170 583026 64226
rect 583094 64170 583150 64226
rect 583218 64170 583274 64226
rect 583342 64170 583398 64226
rect 582970 64046 583026 64102
rect 583094 64046 583150 64102
rect 583218 64046 583274 64102
rect 583342 64046 583398 64102
rect 582970 63922 583026 63978
rect 583094 63922 583150 63978
rect 583218 63922 583274 63978
rect 583342 63922 583398 63978
rect 582970 46294 583026 46350
rect 583094 46294 583150 46350
rect 583218 46294 583274 46350
rect 583342 46294 583398 46350
rect 582970 46170 583026 46226
rect 583094 46170 583150 46226
rect 583218 46170 583274 46226
rect 583342 46170 583398 46226
rect 582970 46046 583026 46102
rect 583094 46046 583150 46102
rect 583218 46046 583274 46102
rect 583342 46046 583398 46102
rect 582970 45922 583026 45978
rect 583094 45922 583150 45978
rect 583218 45922 583274 45978
rect 583342 45922 583398 45978
rect 582970 28294 583026 28350
rect 583094 28294 583150 28350
rect 583218 28294 583274 28350
rect 583342 28294 583398 28350
rect 582970 28170 583026 28226
rect 583094 28170 583150 28226
rect 583218 28170 583274 28226
rect 583342 28170 583398 28226
rect 582970 28046 583026 28102
rect 583094 28046 583150 28102
rect 583218 28046 583274 28102
rect 583342 28046 583398 28102
rect 582970 27922 583026 27978
rect 583094 27922 583150 27978
rect 583218 27922 583274 27978
rect 583342 27922 583398 27978
rect 582970 10294 583026 10350
rect 583094 10294 583150 10350
rect 583218 10294 583274 10350
rect 583342 10294 583398 10350
rect 582970 10170 583026 10226
rect 583094 10170 583150 10226
rect 583218 10170 583274 10226
rect 583342 10170 583398 10226
rect 582970 10046 583026 10102
rect 583094 10046 583150 10102
rect 583218 10046 583274 10102
rect 583342 10046 583398 10102
rect 582970 9922 583026 9978
rect 583094 9922 583150 9978
rect 583218 9922 583274 9978
rect 583342 9922 583398 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 582970 -1176 583026 -1120
rect 583094 -1176 583150 -1120
rect 583218 -1176 583274 -1120
rect 583342 -1176 583398 -1120
rect 582970 -1300 583026 -1244
rect 583094 -1300 583150 -1244
rect 583218 -1300 583274 -1244
rect 583342 -1300 583398 -1244
rect 582970 -1424 583026 -1368
rect 583094 -1424 583150 -1368
rect 583218 -1424 583274 -1368
rect 583342 -1424 583398 -1368
rect 582970 -1548 583026 -1492
rect 583094 -1548 583150 -1492
rect 583218 -1548 583274 -1492
rect 583342 -1548 583398 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 165250 526350
rect 165306 526294 165374 526350
rect 165430 526294 165498 526350
rect 165554 526294 165622 526350
rect 165678 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 255250 526350
rect 255306 526294 255374 526350
rect 255430 526294 255498 526350
rect 255554 526294 255622 526350
rect 255678 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 345250 526350
rect 345306 526294 345374 526350
rect 345430 526294 345498 526350
rect 345554 526294 345622 526350
rect 345678 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 435250 526350
rect 435306 526294 435374 526350
rect 435430 526294 435498 526350
rect 435554 526294 435622 526350
rect 435678 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 525250 526350
rect 525306 526294 525374 526350
rect 525430 526294 525498 526350
rect 525554 526294 525622 526350
rect 525678 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 165250 526226
rect 165306 526170 165374 526226
rect 165430 526170 165498 526226
rect 165554 526170 165622 526226
rect 165678 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 255250 526226
rect 255306 526170 255374 526226
rect 255430 526170 255498 526226
rect 255554 526170 255622 526226
rect 255678 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 345250 526226
rect 345306 526170 345374 526226
rect 345430 526170 345498 526226
rect 345554 526170 345622 526226
rect 345678 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 435250 526226
rect 435306 526170 435374 526226
rect 435430 526170 435498 526226
rect 435554 526170 435622 526226
rect 435678 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 525250 526226
rect 525306 526170 525374 526226
rect 525430 526170 525498 526226
rect 525554 526170 525622 526226
rect 525678 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 165250 526102
rect 165306 526046 165374 526102
rect 165430 526046 165498 526102
rect 165554 526046 165622 526102
rect 165678 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 255250 526102
rect 255306 526046 255374 526102
rect 255430 526046 255498 526102
rect 255554 526046 255622 526102
rect 255678 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 345250 526102
rect 345306 526046 345374 526102
rect 345430 526046 345498 526102
rect 345554 526046 345622 526102
rect 345678 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 435250 526102
rect 435306 526046 435374 526102
rect 435430 526046 435498 526102
rect 435554 526046 435622 526102
rect 435678 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 525250 526102
rect 525306 526046 525374 526102
rect 525430 526046 525498 526102
rect 525554 526046 525622 526102
rect 525678 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 165250 525978
rect 165306 525922 165374 525978
rect 165430 525922 165498 525978
rect 165554 525922 165622 525978
rect 165678 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 255250 525978
rect 255306 525922 255374 525978
rect 255430 525922 255498 525978
rect 255554 525922 255622 525978
rect 255678 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 345250 525978
rect 345306 525922 345374 525978
rect 345430 525922 345498 525978
rect 345554 525922 345622 525978
rect 345678 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 435250 525978
rect 435306 525922 435374 525978
rect 435430 525922 435498 525978
rect 435554 525922 435622 525978
rect 435678 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 525250 525978
rect 525306 525922 525374 525978
rect 525430 525922 525498 525978
rect 525554 525922 525622 525978
rect 525678 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 39878 514350
rect 39934 514294 40002 514350
rect 40058 514294 70598 514350
rect 70654 514294 70722 514350
rect 70778 514294 101318 514350
rect 101374 514294 101442 514350
rect 101498 514294 132038 514350
rect 132094 514294 132162 514350
rect 132218 514294 162758 514350
rect 162814 514294 162882 514350
rect 162938 514294 193478 514350
rect 193534 514294 193602 514350
rect 193658 514294 224198 514350
rect 224254 514294 224322 514350
rect 224378 514294 254918 514350
rect 254974 514294 255042 514350
rect 255098 514294 285638 514350
rect 285694 514294 285762 514350
rect 285818 514294 316358 514350
rect 316414 514294 316482 514350
rect 316538 514294 347078 514350
rect 347134 514294 347202 514350
rect 347258 514294 377798 514350
rect 377854 514294 377922 514350
rect 377978 514294 408518 514350
rect 408574 514294 408642 514350
rect 408698 514294 439238 514350
rect 439294 514294 439362 514350
rect 439418 514294 469958 514350
rect 470014 514294 470082 514350
rect 470138 514294 500678 514350
rect 500734 514294 500802 514350
rect 500858 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 39878 514226
rect 39934 514170 40002 514226
rect 40058 514170 70598 514226
rect 70654 514170 70722 514226
rect 70778 514170 101318 514226
rect 101374 514170 101442 514226
rect 101498 514170 132038 514226
rect 132094 514170 132162 514226
rect 132218 514170 162758 514226
rect 162814 514170 162882 514226
rect 162938 514170 193478 514226
rect 193534 514170 193602 514226
rect 193658 514170 224198 514226
rect 224254 514170 224322 514226
rect 224378 514170 254918 514226
rect 254974 514170 255042 514226
rect 255098 514170 285638 514226
rect 285694 514170 285762 514226
rect 285818 514170 316358 514226
rect 316414 514170 316482 514226
rect 316538 514170 347078 514226
rect 347134 514170 347202 514226
rect 347258 514170 377798 514226
rect 377854 514170 377922 514226
rect 377978 514170 408518 514226
rect 408574 514170 408642 514226
rect 408698 514170 439238 514226
rect 439294 514170 439362 514226
rect 439418 514170 469958 514226
rect 470014 514170 470082 514226
rect 470138 514170 500678 514226
rect 500734 514170 500802 514226
rect 500858 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 39878 514102
rect 39934 514046 40002 514102
rect 40058 514046 70598 514102
rect 70654 514046 70722 514102
rect 70778 514046 101318 514102
rect 101374 514046 101442 514102
rect 101498 514046 132038 514102
rect 132094 514046 132162 514102
rect 132218 514046 162758 514102
rect 162814 514046 162882 514102
rect 162938 514046 193478 514102
rect 193534 514046 193602 514102
rect 193658 514046 224198 514102
rect 224254 514046 224322 514102
rect 224378 514046 254918 514102
rect 254974 514046 255042 514102
rect 255098 514046 285638 514102
rect 285694 514046 285762 514102
rect 285818 514046 316358 514102
rect 316414 514046 316482 514102
rect 316538 514046 347078 514102
rect 347134 514046 347202 514102
rect 347258 514046 377798 514102
rect 377854 514046 377922 514102
rect 377978 514046 408518 514102
rect 408574 514046 408642 514102
rect 408698 514046 439238 514102
rect 439294 514046 439362 514102
rect 439418 514046 469958 514102
rect 470014 514046 470082 514102
rect 470138 514046 500678 514102
rect 500734 514046 500802 514102
rect 500858 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 39878 513978
rect 39934 513922 40002 513978
rect 40058 513922 70598 513978
rect 70654 513922 70722 513978
rect 70778 513922 101318 513978
rect 101374 513922 101442 513978
rect 101498 513922 132038 513978
rect 132094 513922 132162 513978
rect 132218 513922 162758 513978
rect 162814 513922 162882 513978
rect 162938 513922 193478 513978
rect 193534 513922 193602 513978
rect 193658 513922 224198 513978
rect 224254 513922 224322 513978
rect 224378 513922 254918 513978
rect 254974 513922 255042 513978
rect 255098 513922 285638 513978
rect 285694 513922 285762 513978
rect 285818 513922 316358 513978
rect 316414 513922 316482 513978
rect 316538 513922 347078 513978
rect 347134 513922 347202 513978
rect 347258 513922 377798 513978
rect 377854 513922 377922 513978
rect 377978 513922 408518 513978
rect 408574 513922 408642 513978
rect 408698 513922 439238 513978
rect 439294 513922 439362 513978
rect 439418 513922 469958 513978
rect 470014 513922 470082 513978
rect 470138 513922 500678 513978
rect 500734 513922 500802 513978
rect 500858 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 24518 508350
rect 24574 508294 24642 508350
rect 24698 508294 55238 508350
rect 55294 508294 55362 508350
rect 55418 508294 85958 508350
rect 86014 508294 86082 508350
rect 86138 508294 116678 508350
rect 116734 508294 116802 508350
rect 116858 508294 147398 508350
rect 147454 508294 147522 508350
rect 147578 508294 178118 508350
rect 178174 508294 178242 508350
rect 178298 508294 208838 508350
rect 208894 508294 208962 508350
rect 209018 508294 239558 508350
rect 239614 508294 239682 508350
rect 239738 508294 270278 508350
rect 270334 508294 270402 508350
rect 270458 508294 300998 508350
rect 301054 508294 301122 508350
rect 301178 508294 331718 508350
rect 331774 508294 331842 508350
rect 331898 508294 362438 508350
rect 362494 508294 362562 508350
rect 362618 508294 393158 508350
rect 393214 508294 393282 508350
rect 393338 508294 423878 508350
rect 423934 508294 424002 508350
rect 424058 508294 454598 508350
rect 454654 508294 454722 508350
rect 454778 508294 485318 508350
rect 485374 508294 485442 508350
rect 485498 508294 516038 508350
rect 516094 508294 516162 508350
rect 516218 508294 525250 508350
rect 525306 508294 525374 508350
rect 525430 508294 525498 508350
rect 525554 508294 525622 508350
rect 525678 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 24518 508226
rect 24574 508170 24642 508226
rect 24698 508170 55238 508226
rect 55294 508170 55362 508226
rect 55418 508170 85958 508226
rect 86014 508170 86082 508226
rect 86138 508170 116678 508226
rect 116734 508170 116802 508226
rect 116858 508170 147398 508226
rect 147454 508170 147522 508226
rect 147578 508170 178118 508226
rect 178174 508170 178242 508226
rect 178298 508170 208838 508226
rect 208894 508170 208962 508226
rect 209018 508170 239558 508226
rect 239614 508170 239682 508226
rect 239738 508170 270278 508226
rect 270334 508170 270402 508226
rect 270458 508170 300998 508226
rect 301054 508170 301122 508226
rect 301178 508170 331718 508226
rect 331774 508170 331842 508226
rect 331898 508170 362438 508226
rect 362494 508170 362562 508226
rect 362618 508170 393158 508226
rect 393214 508170 393282 508226
rect 393338 508170 423878 508226
rect 423934 508170 424002 508226
rect 424058 508170 454598 508226
rect 454654 508170 454722 508226
rect 454778 508170 485318 508226
rect 485374 508170 485442 508226
rect 485498 508170 516038 508226
rect 516094 508170 516162 508226
rect 516218 508170 525250 508226
rect 525306 508170 525374 508226
rect 525430 508170 525498 508226
rect 525554 508170 525622 508226
rect 525678 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 24518 508102
rect 24574 508046 24642 508102
rect 24698 508046 55238 508102
rect 55294 508046 55362 508102
rect 55418 508046 85958 508102
rect 86014 508046 86082 508102
rect 86138 508046 116678 508102
rect 116734 508046 116802 508102
rect 116858 508046 147398 508102
rect 147454 508046 147522 508102
rect 147578 508046 178118 508102
rect 178174 508046 178242 508102
rect 178298 508046 208838 508102
rect 208894 508046 208962 508102
rect 209018 508046 239558 508102
rect 239614 508046 239682 508102
rect 239738 508046 270278 508102
rect 270334 508046 270402 508102
rect 270458 508046 300998 508102
rect 301054 508046 301122 508102
rect 301178 508046 331718 508102
rect 331774 508046 331842 508102
rect 331898 508046 362438 508102
rect 362494 508046 362562 508102
rect 362618 508046 393158 508102
rect 393214 508046 393282 508102
rect 393338 508046 423878 508102
rect 423934 508046 424002 508102
rect 424058 508046 454598 508102
rect 454654 508046 454722 508102
rect 454778 508046 485318 508102
rect 485374 508046 485442 508102
rect 485498 508046 516038 508102
rect 516094 508046 516162 508102
rect 516218 508046 525250 508102
rect 525306 508046 525374 508102
rect 525430 508046 525498 508102
rect 525554 508046 525622 508102
rect 525678 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 24518 507978
rect 24574 507922 24642 507978
rect 24698 507922 55238 507978
rect 55294 507922 55362 507978
rect 55418 507922 85958 507978
rect 86014 507922 86082 507978
rect 86138 507922 116678 507978
rect 116734 507922 116802 507978
rect 116858 507922 147398 507978
rect 147454 507922 147522 507978
rect 147578 507922 178118 507978
rect 178174 507922 178242 507978
rect 178298 507922 208838 507978
rect 208894 507922 208962 507978
rect 209018 507922 239558 507978
rect 239614 507922 239682 507978
rect 239738 507922 270278 507978
rect 270334 507922 270402 507978
rect 270458 507922 300998 507978
rect 301054 507922 301122 507978
rect 301178 507922 331718 507978
rect 331774 507922 331842 507978
rect 331898 507922 362438 507978
rect 362494 507922 362562 507978
rect 362618 507922 393158 507978
rect 393214 507922 393282 507978
rect 393338 507922 423878 507978
rect 423934 507922 424002 507978
rect 424058 507922 454598 507978
rect 454654 507922 454722 507978
rect 454778 507922 485318 507978
rect 485374 507922 485442 507978
rect 485498 507922 516038 507978
rect 516094 507922 516162 507978
rect 516218 507922 525250 507978
rect 525306 507922 525374 507978
rect 525430 507922 525498 507978
rect 525554 507922 525622 507978
rect 525678 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 39878 496350
rect 39934 496294 40002 496350
rect 40058 496294 70598 496350
rect 70654 496294 70722 496350
rect 70778 496294 101318 496350
rect 101374 496294 101442 496350
rect 101498 496294 132038 496350
rect 132094 496294 132162 496350
rect 132218 496294 162758 496350
rect 162814 496294 162882 496350
rect 162938 496294 193478 496350
rect 193534 496294 193602 496350
rect 193658 496294 224198 496350
rect 224254 496294 224322 496350
rect 224378 496294 254918 496350
rect 254974 496294 255042 496350
rect 255098 496294 285638 496350
rect 285694 496294 285762 496350
rect 285818 496294 316358 496350
rect 316414 496294 316482 496350
rect 316538 496294 347078 496350
rect 347134 496294 347202 496350
rect 347258 496294 377798 496350
rect 377854 496294 377922 496350
rect 377978 496294 408518 496350
rect 408574 496294 408642 496350
rect 408698 496294 439238 496350
rect 439294 496294 439362 496350
rect 439418 496294 469958 496350
rect 470014 496294 470082 496350
rect 470138 496294 500678 496350
rect 500734 496294 500802 496350
rect 500858 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 39878 496226
rect 39934 496170 40002 496226
rect 40058 496170 70598 496226
rect 70654 496170 70722 496226
rect 70778 496170 101318 496226
rect 101374 496170 101442 496226
rect 101498 496170 132038 496226
rect 132094 496170 132162 496226
rect 132218 496170 162758 496226
rect 162814 496170 162882 496226
rect 162938 496170 193478 496226
rect 193534 496170 193602 496226
rect 193658 496170 224198 496226
rect 224254 496170 224322 496226
rect 224378 496170 254918 496226
rect 254974 496170 255042 496226
rect 255098 496170 285638 496226
rect 285694 496170 285762 496226
rect 285818 496170 316358 496226
rect 316414 496170 316482 496226
rect 316538 496170 347078 496226
rect 347134 496170 347202 496226
rect 347258 496170 377798 496226
rect 377854 496170 377922 496226
rect 377978 496170 408518 496226
rect 408574 496170 408642 496226
rect 408698 496170 439238 496226
rect 439294 496170 439362 496226
rect 439418 496170 469958 496226
rect 470014 496170 470082 496226
rect 470138 496170 500678 496226
rect 500734 496170 500802 496226
rect 500858 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 39878 496102
rect 39934 496046 40002 496102
rect 40058 496046 70598 496102
rect 70654 496046 70722 496102
rect 70778 496046 101318 496102
rect 101374 496046 101442 496102
rect 101498 496046 132038 496102
rect 132094 496046 132162 496102
rect 132218 496046 162758 496102
rect 162814 496046 162882 496102
rect 162938 496046 193478 496102
rect 193534 496046 193602 496102
rect 193658 496046 224198 496102
rect 224254 496046 224322 496102
rect 224378 496046 254918 496102
rect 254974 496046 255042 496102
rect 255098 496046 285638 496102
rect 285694 496046 285762 496102
rect 285818 496046 316358 496102
rect 316414 496046 316482 496102
rect 316538 496046 347078 496102
rect 347134 496046 347202 496102
rect 347258 496046 377798 496102
rect 377854 496046 377922 496102
rect 377978 496046 408518 496102
rect 408574 496046 408642 496102
rect 408698 496046 439238 496102
rect 439294 496046 439362 496102
rect 439418 496046 469958 496102
rect 470014 496046 470082 496102
rect 470138 496046 500678 496102
rect 500734 496046 500802 496102
rect 500858 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 39878 495978
rect 39934 495922 40002 495978
rect 40058 495922 70598 495978
rect 70654 495922 70722 495978
rect 70778 495922 101318 495978
rect 101374 495922 101442 495978
rect 101498 495922 132038 495978
rect 132094 495922 132162 495978
rect 132218 495922 162758 495978
rect 162814 495922 162882 495978
rect 162938 495922 193478 495978
rect 193534 495922 193602 495978
rect 193658 495922 224198 495978
rect 224254 495922 224322 495978
rect 224378 495922 254918 495978
rect 254974 495922 255042 495978
rect 255098 495922 285638 495978
rect 285694 495922 285762 495978
rect 285818 495922 316358 495978
rect 316414 495922 316482 495978
rect 316538 495922 347078 495978
rect 347134 495922 347202 495978
rect 347258 495922 377798 495978
rect 377854 495922 377922 495978
rect 377978 495922 408518 495978
rect 408574 495922 408642 495978
rect 408698 495922 439238 495978
rect 439294 495922 439362 495978
rect 439418 495922 469958 495978
rect 470014 495922 470082 495978
rect 470138 495922 500678 495978
rect 500734 495922 500802 495978
rect 500858 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 24518 490350
rect 24574 490294 24642 490350
rect 24698 490294 55238 490350
rect 55294 490294 55362 490350
rect 55418 490294 85958 490350
rect 86014 490294 86082 490350
rect 86138 490294 116678 490350
rect 116734 490294 116802 490350
rect 116858 490294 147398 490350
rect 147454 490294 147522 490350
rect 147578 490294 178118 490350
rect 178174 490294 178242 490350
rect 178298 490294 208838 490350
rect 208894 490294 208962 490350
rect 209018 490294 239558 490350
rect 239614 490294 239682 490350
rect 239738 490294 270278 490350
rect 270334 490294 270402 490350
rect 270458 490294 300998 490350
rect 301054 490294 301122 490350
rect 301178 490294 331718 490350
rect 331774 490294 331842 490350
rect 331898 490294 362438 490350
rect 362494 490294 362562 490350
rect 362618 490294 393158 490350
rect 393214 490294 393282 490350
rect 393338 490294 423878 490350
rect 423934 490294 424002 490350
rect 424058 490294 454598 490350
rect 454654 490294 454722 490350
rect 454778 490294 485318 490350
rect 485374 490294 485442 490350
rect 485498 490294 516038 490350
rect 516094 490294 516162 490350
rect 516218 490294 525250 490350
rect 525306 490294 525374 490350
rect 525430 490294 525498 490350
rect 525554 490294 525622 490350
rect 525678 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 24518 490226
rect 24574 490170 24642 490226
rect 24698 490170 55238 490226
rect 55294 490170 55362 490226
rect 55418 490170 85958 490226
rect 86014 490170 86082 490226
rect 86138 490170 116678 490226
rect 116734 490170 116802 490226
rect 116858 490170 147398 490226
rect 147454 490170 147522 490226
rect 147578 490170 178118 490226
rect 178174 490170 178242 490226
rect 178298 490170 208838 490226
rect 208894 490170 208962 490226
rect 209018 490170 239558 490226
rect 239614 490170 239682 490226
rect 239738 490170 270278 490226
rect 270334 490170 270402 490226
rect 270458 490170 300998 490226
rect 301054 490170 301122 490226
rect 301178 490170 331718 490226
rect 331774 490170 331842 490226
rect 331898 490170 362438 490226
rect 362494 490170 362562 490226
rect 362618 490170 393158 490226
rect 393214 490170 393282 490226
rect 393338 490170 423878 490226
rect 423934 490170 424002 490226
rect 424058 490170 454598 490226
rect 454654 490170 454722 490226
rect 454778 490170 485318 490226
rect 485374 490170 485442 490226
rect 485498 490170 516038 490226
rect 516094 490170 516162 490226
rect 516218 490170 525250 490226
rect 525306 490170 525374 490226
rect 525430 490170 525498 490226
rect 525554 490170 525622 490226
rect 525678 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 24518 490102
rect 24574 490046 24642 490102
rect 24698 490046 55238 490102
rect 55294 490046 55362 490102
rect 55418 490046 85958 490102
rect 86014 490046 86082 490102
rect 86138 490046 116678 490102
rect 116734 490046 116802 490102
rect 116858 490046 147398 490102
rect 147454 490046 147522 490102
rect 147578 490046 178118 490102
rect 178174 490046 178242 490102
rect 178298 490046 208838 490102
rect 208894 490046 208962 490102
rect 209018 490046 239558 490102
rect 239614 490046 239682 490102
rect 239738 490046 270278 490102
rect 270334 490046 270402 490102
rect 270458 490046 300998 490102
rect 301054 490046 301122 490102
rect 301178 490046 331718 490102
rect 331774 490046 331842 490102
rect 331898 490046 362438 490102
rect 362494 490046 362562 490102
rect 362618 490046 393158 490102
rect 393214 490046 393282 490102
rect 393338 490046 423878 490102
rect 423934 490046 424002 490102
rect 424058 490046 454598 490102
rect 454654 490046 454722 490102
rect 454778 490046 485318 490102
rect 485374 490046 485442 490102
rect 485498 490046 516038 490102
rect 516094 490046 516162 490102
rect 516218 490046 525250 490102
rect 525306 490046 525374 490102
rect 525430 490046 525498 490102
rect 525554 490046 525622 490102
rect 525678 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 24518 489978
rect 24574 489922 24642 489978
rect 24698 489922 55238 489978
rect 55294 489922 55362 489978
rect 55418 489922 85958 489978
rect 86014 489922 86082 489978
rect 86138 489922 116678 489978
rect 116734 489922 116802 489978
rect 116858 489922 147398 489978
rect 147454 489922 147522 489978
rect 147578 489922 178118 489978
rect 178174 489922 178242 489978
rect 178298 489922 208838 489978
rect 208894 489922 208962 489978
rect 209018 489922 239558 489978
rect 239614 489922 239682 489978
rect 239738 489922 270278 489978
rect 270334 489922 270402 489978
rect 270458 489922 300998 489978
rect 301054 489922 301122 489978
rect 301178 489922 331718 489978
rect 331774 489922 331842 489978
rect 331898 489922 362438 489978
rect 362494 489922 362562 489978
rect 362618 489922 393158 489978
rect 393214 489922 393282 489978
rect 393338 489922 423878 489978
rect 423934 489922 424002 489978
rect 424058 489922 454598 489978
rect 454654 489922 454722 489978
rect 454778 489922 485318 489978
rect 485374 489922 485442 489978
rect 485498 489922 516038 489978
rect 516094 489922 516162 489978
rect 516218 489922 525250 489978
rect 525306 489922 525374 489978
rect 525430 489922 525498 489978
rect 525554 489922 525622 489978
rect 525678 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 39878 478350
rect 39934 478294 40002 478350
rect 40058 478294 70598 478350
rect 70654 478294 70722 478350
rect 70778 478294 101318 478350
rect 101374 478294 101442 478350
rect 101498 478294 132038 478350
rect 132094 478294 132162 478350
rect 132218 478294 162758 478350
rect 162814 478294 162882 478350
rect 162938 478294 193478 478350
rect 193534 478294 193602 478350
rect 193658 478294 224198 478350
rect 224254 478294 224322 478350
rect 224378 478294 254918 478350
rect 254974 478294 255042 478350
rect 255098 478294 285638 478350
rect 285694 478294 285762 478350
rect 285818 478294 316358 478350
rect 316414 478294 316482 478350
rect 316538 478294 347078 478350
rect 347134 478294 347202 478350
rect 347258 478294 377798 478350
rect 377854 478294 377922 478350
rect 377978 478294 408518 478350
rect 408574 478294 408642 478350
rect 408698 478294 439238 478350
rect 439294 478294 439362 478350
rect 439418 478294 469958 478350
rect 470014 478294 470082 478350
rect 470138 478294 500678 478350
rect 500734 478294 500802 478350
rect 500858 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 39878 478226
rect 39934 478170 40002 478226
rect 40058 478170 70598 478226
rect 70654 478170 70722 478226
rect 70778 478170 101318 478226
rect 101374 478170 101442 478226
rect 101498 478170 132038 478226
rect 132094 478170 132162 478226
rect 132218 478170 162758 478226
rect 162814 478170 162882 478226
rect 162938 478170 193478 478226
rect 193534 478170 193602 478226
rect 193658 478170 224198 478226
rect 224254 478170 224322 478226
rect 224378 478170 254918 478226
rect 254974 478170 255042 478226
rect 255098 478170 285638 478226
rect 285694 478170 285762 478226
rect 285818 478170 316358 478226
rect 316414 478170 316482 478226
rect 316538 478170 347078 478226
rect 347134 478170 347202 478226
rect 347258 478170 377798 478226
rect 377854 478170 377922 478226
rect 377978 478170 408518 478226
rect 408574 478170 408642 478226
rect 408698 478170 439238 478226
rect 439294 478170 439362 478226
rect 439418 478170 469958 478226
rect 470014 478170 470082 478226
rect 470138 478170 500678 478226
rect 500734 478170 500802 478226
rect 500858 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 39878 478102
rect 39934 478046 40002 478102
rect 40058 478046 70598 478102
rect 70654 478046 70722 478102
rect 70778 478046 101318 478102
rect 101374 478046 101442 478102
rect 101498 478046 132038 478102
rect 132094 478046 132162 478102
rect 132218 478046 162758 478102
rect 162814 478046 162882 478102
rect 162938 478046 193478 478102
rect 193534 478046 193602 478102
rect 193658 478046 224198 478102
rect 224254 478046 224322 478102
rect 224378 478046 254918 478102
rect 254974 478046 255042 478102
rect 255098 478046 285638 478102
rect 285694 478046 285762 478102
rect 285818 478046 316358 478102
rect 316414 478046 316482 478102
rect 316538 478046 347078 478102
rect 347134 478046 347202 478102
rect 347258 478046 377798 478102
rect 377854 478046 377922 478102
rect 377978 478046 408518 478102
rect 408574 478046 408642 478102
rect 408698 478046 439238 478102
rect 439294 478046 439362 478102
rect 439418 478046 469958 478102
rect 470014 478046 470082 478102
rect 470138 478046 500678 478102
rect 500734 478046 500802 478102
rect 500858 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 39878 477978
rect 39934 477922 40002 477978
rect 40058 477922 70598 477978
rect 70654 477922 70722 477978
rect 70778 477922 101318 477978
rect 101374 477922 101442 477978
rect 101498 477922 132038 477978
rect 132094 477922 132162 477978
rect 132218 477922 162758 477978
rect 162814 477922 162882 477978
rect 162938 477922 193478 477978
rect 193534 477922 193602 477978
rect 193658 477922 224198 477978
rect 224254 477922 224322 477978
rect 224378 477922 254918 477978
rect 254974 477922 255042 477978
rect 255098 477922 285638 477978
rect 285694 477922 285762 477978
rect 285818 477922 316358 477978
rect 316414 477922 316482 477978
rect 316538 477922 347078 477978
rect 347134 477922 347202 477978
rect 347258 477922 377798 477978
rect 377854 477922 377922 477978
rect 377978 477922 408518 477978
rect 408574 477922 408642 477978
rect 408698 477922 439238 477978
rect 439294 477922 439362 477978
rect 439418 477922 469958 477978
rect 470014 477922 470082 477978
rect 470138 477922 500678 477978
rect 500734 477922 500802 477978
rect 500858 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 24518 472350
rect 24574 472294 24642 472350
rect 24698 472294 55238 472350
rect 55294 472294 55362 472350
rect 55418 472294 85958 472350
rect 86014 472294 86082 472350
rect 86138 472294 116678 472350
rect 116734 472294 116802 472350
rect 116858 472294 147398 472350
rect 147454 472294 147522 472350
rect 147578 472294 178118 472350
rect 178174 472294 178242 472350
rect 178298 472294 208838 472350
rect 208894 472294 208962 472350
rect 209018 472294 239558 472350
rect 239614 472294 239682 472350
rect 239738 472294 270278 472350
rect 270334 472294 270402 472350
rect 270458 472294 300998 472350
rect 301054 472294 301122 472350
rect 301178 472294 331718 472350
rect 331774 472294 331842 472350
rect 331898 472294 362438 472350
rect 362494 472294 362562 472350
rect 362618 472294 393158 472350
rect 393214 472294 393282 472350
rect 393338 472294 423878 472350
rect 423934 472294 424002 472350
rect 424058 472294 454598 472350
rect 454654 472294 454722 472350
rect 454778 472294 485318 472350
rect 485374 472294 485442 472350
rect 485498 472294 516038 472350
rect 516094 472294 516162 472350
rect 516218 472294 525250 472350
rect 525306 472294 525374 472350
rect 525430 472294 525498 472350
rect 525554 472294 525622 472350
rect 525678 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 24518 472226
rect 24574 472170 24642 472226
rect 24698 472170 55238 472226
rect 55294 472170 55362 472226
rect 55418 472170 85958 472226
rect 86014 472170 86082 472226
rect 86138 472170 116678 472226
rect 116734 472170 116802 472226
rect 116858 472170 147398 472226
rect 147454 472170 147522 472226
rect 147578 472170 178118 472226
rect 178174 472170 178242 472226
rect 178298 472170 208838 472226
rect 208894 472170 208962 472226
rect 209018 472170 239558 472226
rect 239614 472170 239682 472226
rect 239738 472170 270278 472226
rect 270334 472170 270402 472226
rect 270458 472170 300998 472226
rect 301054 472170 301122 472226
rect 301178 472170 331718 472226
rect 331774 472170 331842 472226
rect 331898 472170 362438 472226
rect 362494 472170 362562 472226
rect 362618 472170 393158 472226
rect 393214 472170 393282 472226
rect 393338 472170 423878 472226
rect 423934 472170 424002 472226
rect 424058 472170 454598 472226
rect 454654 472170 454722 472226
rect 454778 472170 485318 472226
rect 485374 472170 485442 472226
rect 485498 472170 516038 472226
rect 516094 472170 516162 472226
rect 516218 472170 525250 472226
rect 525306 472170 525374 472226
rect 525430 472170 525498 472226
rect 525554 472170 525622 472226
rect 525678 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 24518 472102
rect 24574 472046 24642 472102
rect 24698 472046 55238 472102
rect 55294 472046 55362 472102
rect 55418 472046 85958 472102
rect 86014 472046 86082 472102
rect 86138 472046 116678 472102
rect 116734 472046 116802 472102
rect 116858 472046 147398 472102
rect 147454 472046 147522 472102
rect 147578 472046 178118 472102
rect 178174 472046 178242 472102
rect 178298 472046 208838 472102
rect 208894 472046 208962 472102
rect 209018 472046 239558 472102
rect 239614 472046 239682 472102
rect 239738 472046 270278 472102
rect 270334 472046 270402 472102
rect 270458 472046 300998 472102
rect 301054 472046 301122 472102
rect 301178 472046 331718 472102
rect 331774 472046 331842 472102
rect 331898 472046 362438 472102
rect 362494 472046 362562 472102
rect 362618 472046 393158 472102
rect 393214 472046 393282 472102
rect 393338 472046 423878 472102
rect 423934 472046 424002 472102
rect 424058 472046 454598 472102
rect 454654 472046 454722 472102
rect 454778 472046 485318 472102
rect 485374 472046 485442 472102
rect 485498 472046 516038 472102
rect 516094 472046 516162 472102
rect 516218 472046 525250 472102
rect 525306 472046 525374 472102
rect 525430 472046 525498 472102
rect 525554 472046 525622 472102
rect 525678 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 24518 471978
rect 24574 471922 24642 471978
rect 24698 471922 55238 471978
rect 55294 471922 55362 471978
rect 55418 471922 85958 471978
rect 86014 471922 86082 471978
rect 86138 471922 116678 471978
rect 116734 471922 116802 471978
rect 116858 471922 147398 471978
rect 147454 471922 147522 471978
rect 147578 471922 178118 471978
rect 178174 471922 178242 471978
rect 178298 471922 208838 471978
rect 208894 471922 208962 471978
rect 209018 471922 239558 471978
rect 239614 471922 239682 471978
rect 239738 471922 270278 471978
rect 270334 471922 270402 471978
rect 270458 471922 300998 471978
rect 301054 471922 301122 471978
rect 301178 471922 331718 471978
rect 331774 471922 331842 471978
rect 331898 471922 362438 471978
rect 362494 471922 362562 471978
rect 362618 471922 393158 471978
rect 393214 471922 393282 471978
rect 393338 471922 423878 471978
rect 423934 471922 424002 471978
rect 424058 471922 454598 471978
rect 454654 471922 454722 471978
rect 454778 471922 485318 471978
rect 485374 471922 485442 471978
rect 485498 471922 516038 471978
rect 516094 471922 516162 471978
rect 516218 471922 525250 471978
rect 525306 471922 525374 471978
rect 525430 471922 525498 471978
rect 525554 471922 525622 471978
rect 525678 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 39878 460350
rect 39934 460294 40002 460350
rect 40058 460294 70598 460350
rect 70654 460294 70722 460350
rect 70778 460294 101318 460350
rect 101374 460294 101442 460350
rect 101498 460294 132038 460350
rect 132094 460294 132162 460350
rect 132218 460294 162758 460350
rect 162814 460294 162882 460350
rect 162938 460294 193478 460350
rect 193534 460294 193602 460350
rect 193658 460294 224198 460350
rect 224254 460294 224322 460350
rect 224378 460294 254918 460350
rect 254974 460294 255042 460350
rect 255098 460294 285638 460350
rect 285694 460294 285762 460350
rect 285818 460294 316358 460350
rect 316414 460294 316482 460350
rect 316538 460294 347078 460350
rect 347134 460294 347202 460350
rect 347258 460294 377798 460350
rect 377854 460294 377922 460350
rect 377978 460294 408518 460350
rect 408574 460294 408642 460350
rect 408698 460294 439238 460350
rect 439294 460294 439362 460350
rect 439418 460294 469958 460350
rect 470014 460294 470082 460350
rect 470138 460294 500678 460350
rect 500734 460294 500802 460350
rect 500858 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 39878 460226
rect 39934 460170 40002 460226
rect 40058 460170 70598 460226
rect 70654 460170 70722 460226
rect 70778 460170 101318 460226
rect 101374 460170 101442 460226
rect 101498 460170 132038 460226
rect 132094 460170 132162 460226
rect 132218 460170 162758 460226
rect 162814 460170 162882 460226
rect 162938 460170 193478 460226
rect 193534 460170 193602 460226
rect 193658 460170 224198 460226
rect 224254 460170 224322 460226
rect 224378 460170 254918 460226
rect 254974 460170 255042 460226
rect 255098 460170 285638 460226
rect 285694 460170 285762 460226
rect 285818 460170 316358 460226
rect 316414 460170 316482 460226
rect 316538 460170 347078 460226
rect 347134 460170 347202 460226
rect 347258 460170 377798 460226
rect 377854 460170 377922 460226
rect 377978 460170 408518 460226
rect 408574 460170 408642 460226
rect 408698 460170 439238 460226
rect 439294 460170 439362 460226
rect 439418 460170 469958 460226
rect 470014 460170 470082 460226
rect 470138 460170 500678 460226
rect 500734 460170 500802 460226
rect 500858 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 39878 460102
rect 39934 460046 40002 460102
rect 40058 460046 70598 460102
rect 70654 460046 70722 460102
rect 70778 460046 101318 460102
rect 101374 460046 101442 460102
rect 101498 460046 132038 460102
rect 132094 460046 132162 460102
rect 132218 460046 162758 460102
rect 162814 460046 162882 460102
rect 162938 460046 193478 460102
rect 193534 460046 193602 460102
rect 193658 460046 224198 460102
rect 224254 460046 224322 460102
rect 224378 460046 254918 460102
rect 254974 460046 255042 460102
rect 255098 460046 285638 460102
rect 285694 460046 285762 460102
rect 285818 460046 316358 460102
rect 316414 460046 316482 460102
rect 316538 460046 347078 460102
rect 347134 460046 347202 460102
rect 347258 460046 377798 460102
rect 377854 460046 377922 460102
rect 377978 460046 408518 460102
rect 408574 460046 408642 460102
rect 408698 460046 439238 460102
rect 439294 460046 439362 460102
rect 439418 460046 469958 460102
rect 470014 460046 470082 460102
rect 470138 460046 500678 460102
rect 500734 460046 500802 460102
rect 500858 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 39878 459978
rect 39934 459922 40002 459978
rect 40058 459922 70598 459978
rect 70654 459922 70722 459978
rect 70778 459922 101318 459978
rect 101374 459922 101442 459978
rect 101498 459922 132038 459978
rect 132094 459922 132162 459978
rect 132218 459922 162758 459978
rect 162814 459922 162882 459978
rect 162938 459922 193478 459978
rect 193534 459922 193602 459978
rect 193658 459922 224198 459978
rect 224254 459922 224322 459978
rect 224378 459922 254918 459978
rect 254974 459922 255042 459978
rect 255098 459922 285638 459978
rect 285694 459922 285762 459978
rect 285818 459922 316358 459978
rect 316414 459922 316482 459978
rect 316538 459922 347078 459978
rect 347134 459922 347202 459978
rect 347258 459922 377798 459978
rect 377854 459922 377922 459978
rect 377978 459922 408518 459978
rect 408574 459922 408642 459978
rect 408698 459922 439238 459978
rect 439294 459922 439362 459978
rect 439418 459922 469958 459978
rect 470014 459922 470082 459978
rect 470138 459922 500678 459978
rect 500734 459922 500802 459978
rect 500858 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 24518 454350
rect 24574 454294 24642 454350
rect 24698 454294 55238 454350
rect 55294 454294 55362 454350
rect 55418 454294 85958 454350
rect 86014 454294 86082 454350
rect 86138 454294 116678 454350
rect 116734 454294 116802 454350
rect 116858 454294 147398 454350
rect 147454 454294 147522 454350
rect 147578 454294 178118 454350
rect 178174 454294 178242 454350
rect 178298 454294 208838 454350
rect 208894 454294 208962 454350
rect 209018 454294 239558 454350
rect 239614 454294 239682 454350
rect 239738 454294 270278 454350
rect 270334 454294 270402 454350
rect 270458 454294 300998 454350
rect 301054 454294 301122 454350
rect 301178 454294 331718 454350
rect 331774 454294 331842 454350
rect 331898 454294 362438 454350
rect 362494 454294 362562 454350
rect 362618 454294 393158 454350
rect 393214 454294 393282 454350
rect 393338 454294 423878 454350
rect 423934 454294 424002 454350
rect 424058 454294 454598 454350
rect 454654 454294 454722 454350
rect 454778 454294 485318 454350
rect 485374 454294 485442 454350
rect 485498 454294 516038 454350
rect 516094 454294 516162 454350
rect 516218 454294 525250 454350
rect 525306 454294 525374 454350
rect 525430 454294 525498 454350
rect 525554 454294 525622 454350
rect 525678 454294 543250 454350
rect 543306 454294 543374 454350
rect 543430 454294 543498 454350
rect 543554 454294 543622 454350
rect 543678 454294 561250 454350
rect 561306 454294 561374 454350
rect 561430 454294 561498 454350
rect 561554 454294 561622 454350
rect 561678 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 24518 454226
rect 24574 454170 24642 454226
rect 24698 454170 55238 454226
rect 55294 454170 55362 454226
rect 55418 454170 85958 454226
rect 86014 454170 86082 454226
rect 86138 454170 116678 454226
rect 116734 454170 116802 454226
rect 116858 454170 147398 454226
rect 147454 454170 147522 454226
rect 147578 454170 178118 454226
rect 178174 454170 178242 454226
rect 178298 454170 208838 454226
rect 208894 454170 208962 454226
rect 209018 454170 239558 454226
rect 239614 454170 239682 454226
rect 239738 454170 270278 454226
rect 270334 454170 270402 454226
rect 270458 454170 300998 454226
rect 301054 454170 301122 454226
rect 301178 454170 331718 454226
rect 331774 454170 331842 454226
rect 331898 454170 362438 454226
rect 362494 454170 362562 454226
rect 362618 454170 393158 454226
rect 393214 454170 393282 454226
rect 393338 454170 423878 454226
rect 423934 454170 424002 454226
rect 424058 454170 454598 454226
rect 454654 454170 454722 454226
rect 454778 454170 485318 454226
rect 485374 454170 485442 454226
rect 485498 454170 516038 454226
rect 516094 454170 516162 454226
rect 516218 454170 525250 454226
rect 525306 454170 525374 454226
rect 525430 454170 525498 454226
rect 525554 454170 525622 454226
rect 525678 454170 543250 454226
rect 543306 454170 543374 454226
rect 543430 454170 543498 454226
rect 543554 454170 543622 454226
rect 543678 454170 561250 454226
rect 561306 454170 561374 454226
rect 561430 454170 561498 454226
rect 561554 454170 561622 454226
rect 561678 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 24518 454102
rect 24574 454046 24642 454102
rect 24698 454046 55238 454102
rect 55294 454046 55362 454102
rect 55418 454046 85958 454102
rect 86014 454046 86082 454102
rect 86138 454046 116678 454102
rect 116734 454046 116802 454102
rect 116858 454046 147398 454102
rect 147454 454046 147522 454102
rect 147578 454046 178118 454102
rect 178174 454046 178242 454102
rect 178298 454046 208838 454102
rect 208894 454046 208962 454102
rect 209018 454046 239558 454102
rect 239614 454046 239682 454102
rect 239738 454046 270278 454102
rect 270334 454046 270402 454102
rect 270458 454046 300998 454102
rect 301054 454046 301122 454102
rect 301178 454046 331718 454102
rect 331774 454046 331842 454102
rect 331898 454046 362438 454102
rect 362494 454046 362562 454102
rect 362618 454046 393158 454102
rect 393214 454046 393282 454102
rect 393338 454046 423878 454102
rect 423934 454046 424002 454102
rect 424058 454046 454598 454102
rect 454654 454046 454722 454102
rect 454778 454046 485318 454102
rect 485374 454046 485442 454102
rect 485498 454046 516038 454102
rect 516094 454046 516162 454102
rect 516218 454046 525250 454102
rect 525306 454046 525374 454102
rect 525430 454046 525498 454102
rect 525554 454046 525622 454102
rect 525678 454046 543250 454102
rect 543306 454046 543374 454102
rect 543430 454046 543498 454102
rect 543554 454046 543622 454102
rect 543678 454046 561250 454102
rect 561306 454046 561374 454102
rect 561430 454046 561498 454102
rect 561554 454046 561622 454102
rect 561678 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 24518 453978
rect 24574 453922 24642 453978
rect 24698 453922 55238 453978
rect 55294 453922 55362 453978
rect 55418 453922 85958 453978
rect 86014 453922 86082 453978
rect 86138 453922 116678 453978
rect 116734 453922 116802 453978
rect 116858 453922 147398 453978
rect 147454 453922 147522 453978
rect 147578 453922 178118 453978
rect 178174 453922 178242 453978
rect 178298 453922 208838 453978
rect 208894 453922 208962 453978
rect 209018 453922 239558 453978
rect 239614 453922 239682 453978
rect 239738 453922 270278 453978
rect 270334 453922 270402 453978
rect 270458 453922 300998 453978
rect 301054 453922 301122 453978
rect 301178 453922 331718 453978
rect 331774 453922 331842 453978
rect 331898 453922 362438 453978
rect 362494 453922 362562 453978
rect 362618 453922 393158 453978
rect 393214 453922 393282 453978
rect 393338 453922 423878 453978
rect 423934 453922 424002 453978
rect 424058 453922 454598 453978
rect 454654 453922 454722 453978
rect 454778 453922 485318 453978
rect 485374 453922 485442 453978
rect 485498 453922 516038 453978
rect 516094 453922 516162 453978
rect 516218 453922 525250 453978
rect 525306 453922 525374 453978
rect 525430 453922 525498 453978
rect 525554 453922 525622 453978
rect 525678 453922 543250 453978
rect 543306 453922 543374 453978
rect 543430 453922 543498 453978
rect 543554 453922 543622 453978
rect 543678 453922 561250 453978
rect 561306 453922 561374 453978
rect 561430 453922 561498 453978
rect 561554 453922 561622 453978
rect 561678 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 39878 442350
rect 39934 442294 40002 442350
rect 40058 442294 70598 442350
rect 70654 442294 70722 442350
rect 70778 442294 101318 442350
rect 101374 442294 101442 442350
rect 101498 442294 132038 442350
rect 132094 442294 132162 442350
rect 132218 442294 162758 442350
rect 162814 442294 162882 442350
rect 162938 442294 193478 442350
rect 193534 442294 193602 442350
rect 193658 442294 224198 442350
rect 224254 442294 224322 442350
rect 224378 442294 254918 442350
rect 254974 442294 255042 442350
rect 255098 442294 285638 442350
rect 285694 442294 285762 442350
rect 285818 442294 316358 442350
rect 316414 442294 316482 442350
rect 316538 442294 347078 442350
rect 347134 442294 347202 442350
rect 347258 442294 377798 442350
rect 377854 442294 377922 442350
rect 377978 442294 408518 442350
rect 408574 442294 408642 442350
rect 408698 442294 439238 442350
rect 439294 442294 439362 442350
rect 439418 442294 469958 442350
rect 470014 442294 470082 442350
rect 470138 442294 500678 442350
rect 500734 442294 500802 442350
rect 500858 442294 528970 442350
rect 529026 442294 529094 442350
rect 529150 442294 529218 442350
rect 529274 442294 529342 442350
rect 529398 442294 546970 442350
rect 547026 442294 547094 442350
rect 547150 442294 547218 442350
rect 547274 442294 547342 442350
rect 547398 442294 564970 442350
rect 565026 442294 565094 442350
rect 565150 442294 565218 442350
rect 565274 442294 565342 442350
rect 565398 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 39878 442226
rect 39934 442170 40002 442226
rect 40058 442170 70598 442226
rect 70654 442170 70722 442226
rect 70778 442170 101318 442226
rect 101374 442170 101442 442226
rect 101498 442170 132038 442226
rect 132094 442170 132162 442226
rect 132218 442170 162758 442226
rect 162814 442170 162882 442226
rect 162938 442170 193478 442226
rect 193534 442170 193602 442226
rect 193658 442170 224198 442226
rect 224254 442170 224322 442226
rect 224378 442170 254918 442226
rect 254974 442170 255042 442226
rect 255098 442170 285638 442226
rect 285694 442170 285762 442226
rect 285818 442170 316358 442226
rect 316414 442170 316482 442226
rect 316538 442170 347078 442226
rect 347134 442170 347202 442226
rect 347258 442170 377798 442226
rect 377854 442170 377922 442226
rect 377978 442170 408518 442226
rect 408574 442170 408642 442226
rect 408698 442170 439238 442226
rect 439294 442170 439362 442226
rect 439418 442170 469958 442226
rect 470014 442170 470082 442226
rect 470138 442170 500678 442226
rect 500734 442170 500802 442226
rect 500858 442170 528970 442226
rect 529026 442170 529094 442226
rect 529150 442170 529218 442226
rect 529274 442170 529342 442226
rect 529398 442170 546970 442226
rect 547026 442170 547094 442226
rect 547150 442170 547218 442226
rect 547274 442170 547342 442226
rect 547398 442170 564970 442226
rect 565026 442170 565094 442226
rect 565150 442170 565218 442226
rect 565274 442170 565342 442226
rect 565398 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 39878 442102
rect 39934 442046 40002 442102
rect 40058 442046 70598 442102
rect 70654 442046 70722 442102
rect 70778 442046 101318 442102
rect 101374 442046 101442 442102
rect 101498 442046 132038 442102
rect 132094 442046 132162 442102
rect 132218 442046 162758 442102
rect 162814 442046 162882 442102
rect 162938 442046 193478 442102
rect 193534 442046 193602 442102
rect 193658 442046 224198 442102
rect 224254 442046 224322 442102
rect 224378 442046 254918 442102
rect 254974 442046 255042 442102
rect 255098 442046 285638 442102
rect 285694 442046 285762 442102
rect 285818 442046 316358 442102
rect 316414 442046 316482 442102
rect 316538 442046 347078 442102
rect 347134 442046 347202 442102
rect 347258 442046 377798 442102
rect 377854 442046 377922 442102
rect 377978 442046 408518 442102
rect 408574 442046 408642 442102
rect 408698 442046 439238 442102
rect 439294 442046 439362 442102
rect 439418 442046 469958 442102
rect 470014 442046 470082 442102
rect 470138 442046 500678 442102
rect 500734 442046 500802 442102
rect 500858 442046 528970 442102
rect 529026 442046 529094 442102
rect 529150 442046 529218 442102
rect 529274 442046 529342 442102
rect 529398 442046 546970 442102
rect 547026 442046 547094 442102
rect 547150 442046 547218 442102
rect 547274 442046 547342 442102
rect 547398 442046 564970 442102
rect 565026 442046 565094 442102
rect 565150 442046 565218 442102
rect 565274 442046 565342 442102
rect 565398 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 39878 441978
rect 39934 441922 40002 441978
rect 40058 441922 70598 441978
rect 70654 441922 70722 441978
rect 70778 441922 101318 441978
rect 101374 441922 101442 441978
rect 101498 441922 132038 441978
rect 132094 441922 132162 441978
rect 132218 441922 162758 441978
rect 162814 441922 162882 441978
rect 162938 441922 193478 441978
rect 193534 441922 193602 441978
rect 193658 441922 224198 441978
rect 224254 441922 224322 441978
rect 224378 441922 254918 441978
rect 254974 441922 255042 441978
rect 255098 441922 285638 441978
rect 285694 441922 285762 441978
rect 285818 441922 316358 441978
rect 316414 441922 316482 441978
rect 316538 441922 347078 441978
rect 347134 441922 347202 441978
rect 347258 441922 377798 441978
rect 377854 441922 377922 441978
rect 377978 441922 408518 441978
rect 408574 441922 408642 441978
rect 408698 441922 439238 441978
rect 439294 441922 439362 441978
rect 439418 441922 469958 441978
rect 470014 441922 470082 441978
rect 470138 441922 500678 441978
rect 500734 441922 500802 441978
rect 500858 441922 528970 441978
rect 529026 441922 529094 441978
rect 529150 441922 529218 441978
rect 529274 441922 529342 441978
rect 529398 441922 546970 441978
rect 547026 441922 547094 441978
rect 547150 441922 547218 441978
rect 547274 441922 547342 441978
rect 547398 441922 564970 441978
rect 565026 441922 565094 441978
rect 565150 441922 565218 441978
rect 565274 441922 565342 441978
rect 565398 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 24518 436350
rect 24574 436294 24642 436350
rect 24698 436294 55238 436350
rect 55294 436294 55362 436350
rect 55418 436294 85958 436350
rect 86014 436294 86082 436350
rect 86138 436294 116678 436350
rect 116734 436294 116802 436350
rect 116858 436294 147398 436350
rect 147454 436294 147522 436350
rect 147578 436294 178118 436350
rect 178174 436294 178242 436350
rect 178298 436294 208838 436350
rect 208894 436294 208962 436350
rect 209018 436294 239558 436350
rect 239614 436294 239682 436350
rect 239738 436294 270278 436350
rect 270334 436294 270402 436350
rect 270458 436294 300998 436350
rect 301054 436294 301122 436350
rect 301178 436294 331718 436350
rect 331774 436294 331842 436350
rect 331898 436294 362438 436350
rect 362494 436294 362562 436350
rect 362618 436294 393158 436350
rect 393214 436294 393282 436350
rect 393338 436294 423878 436350
rect 423934 436294 424002 436350
rect 424058 436294 454598 436350
rect 454654 436294 454722 436350
rect 454778 436294 485318 436350
rect 485374 436294 485442 436350
rect 485498 436294 516038 436350
rect 516094 436294 516162 436350
rect 516218 436294 525250 436350
rect 525306 436294 525374 436350
rect 525430 436294 525498 436350
rect 525554 436294 525622 436350
rect 525678 436294 543250 436350
rect 543306 436294 543374 436350
rect 543430 436294 543498 436350
rect 543554 436294 543622 436350
rect 543678 436294 561250 436350
rect 561306 436294 561374 436350
rect 561430 436294 561498 436350
rect 561554 436294 561622 436350
rect 561678 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 24518 436226
rect 24574 436170 24642 436226
rect 24698 436170 55238 436226
rect 55294 436170 55362 436226
rect 55418 436170 85958 436226
rect 86014 436170 86082 436226
rect 86138 436170 116678 436226
rect 116734 436170 116802 436226
rect 116858 436170 147398 436226
rect 147454 436170 147522 436226
rect 147578 436170 178118 436226
rect 178174 436170 178242 436226
rect 178298 436170 208838 436226
rect 208894 436170 208962 436226
rect 209018 436170 239558 436226
rect 239614 436170 239682 436226
rect 239738 436170 270278 436226
rect 270334 436170 270402 436226
rect 270458 436170 300998 436226
rect 301054 436170 301122 436226
rect 301178 436170 331718 436226
rect 331774 436170 331842 436226
rect 331898 436170 362438 436226
rect 362494 436170 362562 436226
rect 362618 436170 393158 436226
rect 393214 436170 393282 436226
rect 393338 436170 423878 436226
rect 423934 436170 424002 436226
rect 424058 436170 454598 436226
rect 454654 436170 454722 436226
rect 454778 436170 485318 436226
rect 485374 436170 485442 436226
rect 485498 436170 516038 436226
rect 516094 436170 516162 436226
rect 516218 436170 525250 436226
rect 525306 436170 525374 436226
rect 525430 436170 525498 436226
rect 525554 436170 525622 436226
rect 525678 436170 543250 436226
rect 543306 436170 543374 436226
rect 543430 436170 543498 436226
rect 543554 436170 543622 436226
rect 543678 436170 561250 436226
rect 561306 436170 561374 436226
rect 561430 436170 561498 436226
rect 561554 436170 561622 436226
rect 561678 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 24518 436102
rect 24574 436046 24642 436102
rect 24698 436046 55238 436102
rect 55294 436046 55362 436102
rect 55418 436046 85958 436102
rect 86014 436046 86082 436102
rect 86138 436046 116678 436102
rect 116734 436046 116802 436102
rect 116858 436046 147398 436102
rect 147454 436046 147522 436102
rect 147578 436046 178118 436102
rect 178174 436046 178242 436102
rect 178298 436046 208838 436102
rect 208894 436046 208962 436102
rect 209018 436046 239558 436102
rect 239614 436046 239682 436102
rect 239738 436046 270278 436102
rect 270334 436046 270402 436102
rect 270458 436046 300998 436102
rect 301054 436046 301122 436102
rect 301178 436046 331718 436102
rect 331774 436046 331842 436102
rect 331898 436046 362438 436102
rect 362494 436046 362562 436102
rect 362618 436046 393158 436102
rect 393214 436046 393282 436102
rect 393338 436046 423878 436102
rect 423934 436046 424002 436102
rect 424058 436046 454598 436102
rect 454654 436046 454722 436102
rect 454778 436046 485318 436102
rect 485374 436046 485442 436102
rect 485498 436046 516038 436102
rect 516094 436046 516162 436102
rect 516218 436046 525250 436102
rect 525306 436046 525374 436102
rect 525430 436046 525498 436102
rect 525554 436046 525622 436102
rect 525678 436046 543250 436102
rect 543306 436046 543374 436102
rect 543430 436046 543498 436102
rect 543554 436046 543622 436102
rect 543678 436046 561250 436102
rect 561306 436046 561374 436102
rect 561430 436046 561498 436102
rect 561554 436046 561622 436102
rect 561678 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 24518 435978
rect 24574 435922 24642 435978
rect 24698 435922 55238 435978
rect 55294 435922 55362 435978
rect 55418 435922 85958 435978
rect 86014 435922 86082 435978
rect 86138 435922 116678 435978
rect 116734 435922 116802 435978
rect 116858 435922 147398 435978
rect 147454 435922 147522 435978
rect 147578 435922 178118 435978
rect 178174 435922 178242 435978
rect 178298 435922 208838 435978
rect 208894 435922 208962 435978
rect 209018 435922 239558 435978
rect 239614 435922 239682 435978
rect 239738 435922 270278 435978
rect 270334 435922 270402 435978
rect 270458 435922 300998 435978
rect 301054 435922 301122 435978
rect 301178 435922 331718 435978
rect 331774 435922 331842 435978
rect 331898 435922 362438 435978
rect 362494 435922 362562 435978
rect 362618 435922 393158 435978
rect 393214 435922 393282 435978
rect 393338 435922 423878 435978
rect 423934 435922 424002 435978
rect 424058 435922 454598 435978
rect 454654 435922 454722 435978
rect 454778 435922 485318 435978
rect 485374 435922 485442 435978
rect 485498 435922 516038 435978
rect 516094 435922 516162 435978
rect 516218 435922 525250 435978
rect 525306 435922 525374 435978
rect 525430 435922 525498 435978
rect 525554 435922 525622 435978
rect 525678 435922 543250 435978
rect 543306 435922 543374 435978
rect 543430 435922 543498 435978
rect 543554 435922 543622 435978
rect 543678 435922 561250 435978
rect 561306 435922 561374 435978
rect 561430 435922 561498 435978
rect 561554 435922 561622 435978
rect 561678 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 39878 424350
rect 39934 424294 40002 424350
rect 40058 424294 70598 424350
rect 70654 424294 70722 424350
rect 70778 424294 101318 424350
rect 101374 424294 101442 424350
rect 101498 424294 132038 424350
rect 132094 424294 132162 424350
rect 132218 424294 162758 424350
rect 162814 424294 162882 424350
rect 162938 424294 193478 424350
rect 193534 424294 193602 424350
rect 193658 424294 224198 424350
rect 224254 424294 224322 424350
rect 224378 424294 254918 424350
rect 254974 424294 255042 424350
rect 255098 424294 285638 424350
rect 285694 424294 285762 424350
rect 285818 424294 316358 424350
rect 316414 424294 316482 424350
rect 316538 424294 347078 424350
rect 347134 424294 347202 424350
rect 347258 424294 377798 424350
rect 377854 424294 377922 424350
rect 377978 424294 408518 424350
rect 408574 424294 408642 424350
rect 408698 424294 439238 424350
rect 439294 424294 439362 424350
rect 439418 424294 469958 424350
rect 470014 424294 470082 424350
rect 470138 424294 500678 424350
rect 500734 424294 500802 424350
rect 500858 424294 528970 424350
rect 529026 424294 529094 424350
rect 529150 424294 529218 424350
rect 529274 424294 529342 424350
rect 529398 424294 546970 424350
rect 547026 424294 547094 424350
rect 547150 424294 547218 424350
rect 547274 424294 547342 424350
rect 547398 424294 564970 424350
rect 565026 424294 565094 424350
rect 565150 424294 565218 424350
rect 565274 424294 565342 424350
rect 565398 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 39878 424226
rect 39934 424170 40002 424226
rect 40058 424170 70598 424226
rect 70654 424170 70722 424226
rect 70778 424170 101318 424226
rect 101374 424170 101442 424226
rect 101498 424170 132038 424226
rect 132094 424170 132162 424226
rect 132218 424170 162758 424226
rect 162814 424170 162882 424226
rect 162938 424170 193478 424226
rect 193534 424170 193602 424226
rect 193658 424170 224198 424226
rect 224254 424170 224322 424226
rect 224378 424170 254918 424226
rect 254974 424170 255042 424226
rect 255098 424170 285638 424226
rect 285694 424170 285762 424226
rect 285818 424170 316358 424226
rect 316414 424170 316482 424226
rect 316538 424170 347078 424226
rect 347134 424170 347202 424226
rect 347258 424170 377798 424226
rect 377854 424170 377922 424226
rect 377978 424170 408518 424226
rect 408574 424170 408642 424226
rect 408698 424170 439238 424226
rect 439294 424170 439362 424226
rect 439418 424170 469958 424226
rect 470014 424170 470082 424226
rect 470138 424170 500678 424226
rect 500734 424170 500802 424226
rect 500858 424170 528970 424226
rect 529026 424170 529094 424226
rect 529150 424170 529218 424226
rect 529274 424170 529342 424226
rect 529398 424170 546970 424226
rect 547026 424170 547094 424226
rect 547150 424170 547218 424226
rect 547274 424170 547342 424226
rect 547398 424170 564970 424226
rect 565026 424170 565094 424226
rect 565150 424170 565218 424226
rect 565274 424170 565342 424226
rect 565398 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 39878 424102
rect 39934 424046 40002 424102
rect 40058 424046 70598 424102
rect 70654 424046 70722 424102
rect 70778 424046 101318 424102
rect 101374 424046 101442 424102
rect 101498 424046 132038 424102
rect 132094 424046 132162 424102
rect 132218 424046 162758 424102
rect 162814 424046 162882 424102
rect 162938 424046 193478 424102
rect 193534 424046 193602 424102
rect 193658 424046 224198 424102
rect 224254 424046 224322 424102
rect 224378 424046 254918 424102
rect 254974 424046 255042 424102
rect 255098 424046 285638 424102
rect 285694 424046 285762 424102
rect 285818 424046 316358 424102
rect 316414 424046 316482 424102
rect 316538 424046 347078 424102
rect 347134 424046 347202 424102
rect 347258 424046 377798 424102
rect 377854 424046 377922 424102
rect 377978 424046 408518 424102
rect 408574 424046 408642 424102
rect 408698 424046 439238 424102
rect 439294 424046 439362 424102
rect 439418 424046 469958 424102
rect 470014 424046 470082 424102
rect 470138 424046 500678 424102
rect 500734 424046 500802 424102
rect 500858 424046 528970 424102
rect 529026 424046 529094 424102
rect 529150 424046 529218 424102
rect 529274 424046 529342 424102
rect 529398 424046 546970 424102
rect 547026 424046 547094 424102
rect 547150 424046 547218 424102
rect 547274 424046 547342 424102
rect 547398 424046 564970 424102
rect 565026 424046 565094 424102
rect 565150 424046 565218 424102
rect 565274 424046 565342 424102
rect 565398 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 39878 423978
rect 39934 423922 40002 423978
rect 40058 423922 70598 423978
rect 70654 423922 70722 423978
rect 70778 423922 101318 423978
rect 101374 423922 101442 423978
rect 101498 423922 132038 423978
rect 132094 423922 132162 423978
rect 132218 423922 162758 423978
rect 162814 423922 162882 423978
rect 162938 423922 193478 423978
rect 193534 423922 193602 423978
rect 193658 423922 224198 423978
rect 224254 423922 224322 423978
rect 224378 423922 254918 423978
rect 254974 423922 255042 423978
rect 255098 423922 285638 423978
rect 285694 423922 285762 423978
rect 285818 423922 316358 423978
rect 316414 423922 316482 423978
rect 316538 423922 347078 423978
rect 347134 423922 347202 423978
rect 347258 423922 377798 423978
rect 377854 423922 377922 423978
rect 377978 423922 408518 423978
rect 408574 423922 408642 423978
rect 408698 423922 439238 423978
rect 439294 423922 439362 423978
rect 439418 423922 469958 423978
rect 470014 423922 470082 423978
rect 470138 423922 500678 423978
rect 500734 423922 500802 423978
rect 500858 423922 528970 423978
rect 529026 423922 529094 423978
rect 529150 423922 529218 423978
rect 529274 423922 529342 423978
rect 529398 423922 546970 423978
rect 547026 423922 547094 423978
rect 547150 423922 547218 423978
rect 547274 423922 547342 423978
rect 547398 423922 564970 423978
rect 565026 423922 565094 423978
rect 565150 423922 565218 423978
rect 565274 423922 565342 423978
rect 565398 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 24518 418350
rect 24574 418294 24642 418350
rect 24698 418294 55238 418350
rect 55294 418294 55362 418350
rect 55418 418294 85958 418350
rect 86014 418294 86082 418350
rect 86138 418294 116678 418350
rect 116734 418294 116802 418350
rect 116858 418294 147398 418350
rect 147454 418294 147522 418350
rect 147578 418294 178118 418350
rect 178174 418294 178242 418350
rect 178298 418294 208838 418350
rect 208894 418294 208962 418350
rect 209018 418294 239558 418350
rect 239614 418294 239682 418350
rect 239738 418294 270278 418350
rect 270334 418294 270402 418350
rect 270458 418294 300998 418350
rect 301054 418294 301122 418350
rect 301178 418294 331718 418350
rect 331774 418294 331842 418350
rect 331898 418294 362438 418350
rect 362494 418294 362562 418350
rect 362618 418294 393158 418350
rect 393214 418294 393282 418350
rect 393338 418294 423878 418350
rect 423934 418294 424002 418350
rect 424058 418294 454598 418350
rect 454654 418294 454722 418350
rect 454778 418294 485318 418350
rect 485374 418294 485442 418350
rect 485498 418294 516038 418350
rect 516094 418294 516162 418350
rect 516218 418294 525250 418350
rect 525306 418294 525374 418350
rect 525430 418294 525498 418350
rect 525554 418294 525622 418350
rect 525678 418294 543250 418350
rect 543306 418294 543374 418350
rect 543430 418294 543498 418350
rect 543554 418294 543622 418350
rect 543678 418294 561250 418350
rect 561306 418294 561374 418350
rect 561430 418294 561498 418350
rect 561554 418294 561622 418350
rect 561678 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 24518 418226
rect 24574 418170 24642 418226
rect 24698 418170 55238 418226
rect 55294 418170 55362 418226
rect 55418 418170 85958 418226
rect 86014 418170 86082 418226
rect 86138 418170 116678 418226
rect 116734 418170 116802 418226
rect 116858 418170 147398 418226
rect 147454 418170 147522 418226
rect 147578 418170 178118 418226
rect 178174 418170 178242 418226
rect 178298 418170 208838 418226
rect 208894 418170 208962 418226
rect 209018 418170 239558 418226
rect 239614 418170 239682 418226
rect 239738 418170 270278 418226
rect 270334 418170 270402 418226
rect 270458 418170 300998 418226
rect 301054 418170 301122 418226
rect 301178 418170 331718 418226
rect 331774 418170 331842 418226
rect 331898 418170 362438 418226
rect 362494 418170 362562 418226
rect 362618 418170 393158 418226
rect 393214 418170 393282 418226
rect 393338 418170 423878 418226
rect 423934 418170 424002 418226
rect 424058 418170 454598 418226
rect 454654 418170 454722 418226
rect 454778 418170 485318 418226
rect 485374 418170 485442 418226
rect 485498 418170 516038 418226
rect 516094 418170 516162 418226
rect 516218 418170 525250 418226
rect 525306 418170 525374 418226
rect 525430 418170 525498 418226
rect 525554 418170 525622 418226
rect 525678 418170 543250 418226
rect 543306 418170 543374 418226
rect 543430 418170 543498 418226
rect 543554 418170 543622 418226
rect 543678 418170 561250 418226
rect 561306 418170 561374 418226
rect 561430 418170 561498 418226
rect 561554 418170 561622 418226
rect 561678 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 24518 418102
rect 24574 418046 24642 418102
rect 24698 418046 55238 418102
rect 55294 418046 55362 418102
rect 55418 418046 85958 418102
rect 86014 418046 86082 418102
rect 86138 418046 116678 418102
rect 116734 418046 116802 418102
rect 116858 418046 147398 418102
rect 147454 418046 147522 418102
rect 147578 418046 178118 418102
rect 178174 418046 178242 418102
rect 178298 418046 208838 418102
rect 208894 418046 208962 418102
rect 209018 418046 239558 418102
rect 239614 418046 239682 418102
rect 239738 418046 270278 418102
rect 270334 418046 270402 418102
rect 270458 418046 300998 418102
rect 301054 418046 301122 418102
rect 301178 418046 331718 418102
rect 331774 418046 331842 418102
rect 331898 418046 362438 418102
rect 362494 418046 362562 418102
rect 362618 418046 393158 418102
rect 393214 418046 393282 418102
rect 393338 418046 423878 418102
rect 423934 418046 424002 418102
rect 424058 418046 454598 418102
rect 454654 418046 454722 418102
rect 454778 418046 485318 418102
rect 485374 418046 485442 418102
rect 485498 418046 516038 418102
rect 516094 418046 516162 418102
rect 516218 418046 525250 418102
rect 525306 418046 525374 418102
rect 525430 418046 525498 418102
rect 525554 418046 525622 418102
rect 525678 418046 543250 418102
rect 543306 418046 543374 418102
rect 543430 418046 543498 418102
rect 543554 418046 543622 418102
rect 543678 418046 561250 418102
rect 561306 418046 561374 418102
rect 561430 418046 561498 418102
rect 561554 418046 561622 418102
rect 561678 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 24518 417978
rect 24574 417922 24642 417978
rect 24698 417922 55238 417978
rect 55294 417922 55362 417978
rect 55418 417922 85958 417978
rect 86014 417922 86082 417978
rect 86138 417922 116678 417978
rect 116734 417922 116802 417978
rect 116858 417922 147398 417978
rect 147454 417922 147522 417978
rect 147578 417922 178118 417978
rect 178174 417922 178242 417978
rect 178298 417922 208838 417978
rect 208894 417922 208962 417978
rect 209018 417922 239558 417978
rect 239614 417922 239682 417978
rect 239738 417922 270278 417978
rect 270334 417922 270402 417978
rect 270458 417922 300998 417978
rect 301054 417922 301122 417978
rect 301178 417922 331718 417978
rect 331774 417922 331842 417978
rect 331898 417922 362438 417978
rect 362494 417922 362562 417978
rect 362618 417922 393158 417978
rect 393214 417922 393282 417978
rect 393338 417922 423878 417978
rect 423934 417922 424002 417978
rect 424058 417922 454598 417978
rect 454654 417922 454722 417978
rect 454778 417922 485318 417978
rect 485374 417922 485442 417978
rect 485498 417922 516038 417978
rect 516094 417922 516162 417978
rect 516218 417922 525250 417978
rect 525306 417922 525374 417978
rect 525430 417922 525498 417978
rect 525554 417922 525622 417978
rect 525678 417922 543250 417978
rect 543306 417922 543374 417978
rect 543430 417922 543498 417978
rect 543554 417922 543622 417978
rect 543678 417922 561250 417978
rect 561306 417922 561374 417978
rect 561430 417922 561498 417978
rect 561554 417922 561622 417978
rect 561678 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 39878 406350
rect 39934 406294 40002 406350
rect 40058 406294 70598 406350
rect 70654 406294 70722 406350
rect 70778 406294 101318 406350
rect 101374 406294 101442 406350
rect 101498 406294 132038 406350
rect 132094 406294 132162 406350
rect 132218 406294 162758 406350
rect 162814 406294 162882 406350
rect 162938 406294 193478 406350
rect 193534 406294 193602 406350
rect 193658 406294 224198 406350
rect 224254 406294 224322 406350
rect 224378 406294 254918 406350
rect 254974 406294 255042 406350
rect 255098 406294 285638 406350
rect 285694 406294 285762 406350
rect 285818 406294 316358 406350
rect 316414 406294 316482 406350
rect 316538 406294 347078 406350
rect 347134 406294 347202 406350
rect 347258 406294 377798 406350
rect 377854 406294 377922 406350
rect 377978 406294 408518 406350
rect 408574 406294 408642 406350
rect 408698 406294 439238 406350
rect 439294 406294 439362 406350
rect 439418 406294 469958 406350
rect 470014 406294 470082 406350
rect 470138 406294 500678 406350
rect 500734 406294 500802 406350
rect 500858 406294 528970 406350
rect 529026 406294 529094 406350
rect 529150 406294 529218 406350
rect 529274 406294 529342 406350
rect 529398 406294 546970 406350
rect 547026 406294 547094 406350
rect 547150 406294 547218 406350
rect 547274 406294 547342 406350
rect 547398 406294 564970 406350
rect 565026 406294 565094 406350
rect 565150 406294 565218 406350
rect 565274 406294 565342 406350
rect 565398 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 39878 406226
rect 39934 406170 40002 406226
rect 40058 406170 70598 406226
rect 70654 406170 70722 406226
rect 70778 406170 101318 406226
rect 101374 406170 101442 406226
rect 101498 406170 132038 406226
rect 132094 406170 132162 406226
rect 132218 406170 162758 406226
rect 162814 406170 162882 406226
rect 162938 406170 193478 406226
rect 193534 406170 193602 406226
rect 193658 406170 224198 406226
rect 224254 406170 224322 406226
rect 224378 406170 254918 406226
rect 254974 406170 255042 406226
rect 255098 406170 285638 406226
rect 285694 406170 285762 406226
rect 285818 406170 316358 406226
rect 316414 406170 316482 406226
rect 316538 406170 347078 406226
rect 347134 406170 347202 406226
rect 347258 406170 377798 406226
rect 377854 406170 377922 406226
rect 377978 406170 408518 406226
rect 408574 406170 408642 406226
rect 408698 406170 439238 406226
rect 439294 406170 439362 406226
rect 439418 406170 469958 406226
rect 470014 406170 470082 406226
rect 470138 406170 500678 406226
rect 500734 406170 500802 406226
rect 500858 406170 528970 406226
rect 529026 406170 529094 406226
rect 529150 406170 529218 406226
rect 529274 406170 529342 406226
rect 529398 406170 546970 406226
rect 547026 406170 547094 406226
rect 547150 406170 547218 406226
rect 547274 406170 547342 406226
rect 547398 406170 564970 406226
rect 565026 406170 565094 406226
rect 565150 406170 565218 406226
rect 565274 406170 565342 406226
rect 565398 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 39878 406102
rect 39934 406046 40002 406102
rect 40058 406046 70598 406102
rect 70654 406046 70722 406102
rect 70778 406046 101318 406102
rect 101374 406046 101442 406102
rect 101498 406046 132038 406102
rect 132094 406046 132162 406102
rect 132218 406046 162758 406102
rect 162814 406046 162882 406102
rect 162938 406046 193478 406102
rect 193534 406046 193602 406102
rect 193658 406046 224198 406102
rect 224254 406046 224322 406102
rect 224378 406046 254918 406102
rect 254974 406046 255042 406102
rect 255098 406046 285638 406102
rect 285694 406046 285762 406102
rect 285818 406046 316358 406102
rect 316414 406046 316482 406102
rect 316538 406046 347078 406102
rect 347134 406046 347202 406102
rect 347258 406046 377798 406102
rect 377854 406046 377922 406102
rect 377978 406046 408518 406102
rect 408574 406046 408642 406102
rect 408698 406046 439238 406102
rect 439294 406046 439362 406102
rect 439418 406046 469958 406102
rect 470014 406046 470082 406102
rect 470138 406046 500678 406102
rect 500734 406046 500802 406102
rect 500858 406046 528970 406102
rect 529026 406046 529094 406102
rect 529150 406046 529218 406102
rect 529274 406046 529342 406102
rect 529398 406046 546970 406102
rect 547026 406046 547094 406102
rect 547150 406046 547218 406102
rect 547274 406046 547342 406102
rect 547398 406046 564970 406102
rect 565026 406046 565094 406102
rect 565150 406046 565218 406102
rect 565274 406046 565342 406102
rect 565398 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 39878 405978
rect 39934 405922 40002 405978
rect 40058 405922 70598 405978
rect 70654 405922 70722 405978
rect 70778 405922 101318 405978
rect 101374 405922 101442 405978
rect 101498 405922 132038 405978
rect 132094 405922 132162 405978
rect 132218 405922 162758 405978
rect 162814 405922 162882 405978
rect 162938 405922 193478 405978
rect 193534 405922 193602 405978
rect 193658 405922 224198 405978
rect 224254 405922 224322 405978
rect 224378 405922 254918 405978
rect 254974 405922 255042 405978
rect 255098 405922 285638 405978
rect 285694 405922 285762 405978
rect 285818 405922 316358 405978
rect 316414 405922 316482 405978
rect 316538 405922 347078 405978
rect 347134 405922 347202 405978
rect 347258 405922 377798 405978
rect 377854 405922 377922 405978
rect 377978 405922 408518 405978
rect 408574 405922 408642 405978
rect 408698 405922 439238 405978
rect 439294 405922 439362 405978
rect 439418 405922 469958 405978
rect 470014 405922 470082 405978
rect 470138 405922 500678 405978
rect 500734 405922 500802 405978
rect 500858 405922 528970 405978
rect 529026 405922 529094 405978
rect 529150 405922 529218 405978
rect 529274 405922 529342 405978
rect 529398 405922 546970 405978
rect 547026 405922 547094 405978
rect 547150 405922 547218 405978
rect 547274 405922 547342 405978
rect 547398 405922 564970 405978
rect 565026 405922 565094 405978
rect 565150 405922 565218 405978
rect 565274 405922 565342 405978
rect 565398 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 24518 400350
rect 24574 400294 24642 400350
rect 24698 400294 55238 400350
rect 55294 400294 55362 400350
rect 55418 400294 85958 400350
rect 86014 400294 86082 400350
rect 86138 400294 116678 400350
rect 116734 400294 116802 400350
rect 116858 400294 147398 400350
rect 147454 400294 147522 400350
rect 147578 400294 178118 400350
rect 178174 400294 178242 400350
rect 178298 400294 208838 400350
rect 208894 400294 208962 400350
rect 209018 400294 239558 400350
rect 239614 400294 239682 400350
rect 239738 400294 270278 400350
rect 270334 400294 270402 400350
rect 270458 400294 300998 400350
rect 301054 400294 301122 400350
rect 301178 400294 331718 400350
rect 331774 400294 331842 400350
rect 331898 400294 362438 400350
rect 362494 400294 362562 400350
rect 362618 400294 393158 400350
rect 393214 400294 393282 400350
rect 393338 400294 423878 400350
rect 423934 400294 424002 400350
rect 424058 400294 454598 400350
rect 454654 400294 454722 400350
rect 454778 400294 485318 400350
rect 485374 400294 485442 400350
rect 485498 400294 516038 400350
rect 516094 400294 516162 400350
rect 516218 400294 525250 400350
rect 525306 400294 525374 400350
rect 525430 400294 525498 400350
rect 525554 400294 525622 400350
rect 525678 400294 543250 400350
rect 543306 400294 543374 400350
rect 543430 400294 543498 400350
rect 543554 400294 543622 400350
rect 543678 400294 561250 400350
rect 561306 400294 561374 400350
rect 561430 400294 561498 400350
rect 561554 400294 561622 400350
rect 561678 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 24518 400226
rect 24574 400170 24642 400226
rect 24698 400170 55238 400226
rect 55294 400170 55362 400226
rect 55418 400170 85958 400226
rect 86014 400170 86082 400226
rect 86138 400170 116678 400226
rect 116734 400170 116802 400226
rect 116858 400170 147398 400226
rect 147454 400170 147522 400226
rect 147578 400170 178118 400226
rect 178174 400170 178242 400226
rect 178298 400170 208838 400226
rect 208894 400170 208962 400226
rect 209018 400170 239558 400226
rect 239614 400170 239682 400226
rect 239738 400170 270278 400226
rect 270334 400170 270402 400226
rect 270458 400170 300998 400226
rect 301054 400170 301122 400226
rect 301178 400170 331718 400226
rect 331774 400170 331842 400226
rect 331898 400170 362438 400226
rect 362494 400170 362562 400226
rect 362618 400170 393158 400226
rect 393214 400170 393282 400226
rect 393338 400170 423878 400226
rect 423934 400170 424002 400226
rect 424058 400170 454598 400226
rect 454654 400170 454722 400226
rect 454778 400170 485318 400226
rect 485374 400170 485442 400226
rect 485498 400170 516038 400226
rect 516094 400170 516162 400226
rect 516218 400170 525250 400226
rect 525306 400170 525374 400226
rect 525430 400170 525498 400226
rect 525554 400170 525622 400226
rect 525678 400170 543250 400226
rect 543306 400170 543374 400226
rect 543430 400170 543498 400226
rect 543554 400170 543622 400226
rect 543678 400170 561250 400226
rect 561306 400170 561374 400226
rect 561430 400170 561498 400226
rect 561554 400170 561622 400226
rect 561678 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 24518 400102
rect 24574 400046 24642 400102
rect 24698 400046 55238 400102
rect 55294 400046 55362 400102
rect 55418 400046 85958 400102
rect 86014 400046 86082 400102
rect 86138 400046 116678 400102
rect 116734 400046 116802 400102
rect 116858 400046 147398 400102
rect 147454 400046 147522 400102
rect 147578 400046 178118 400102
rect 178174 400046 178242 400102
rect 178298 400046 208838 400102
rect 208894 400046 208962 400102
rect 209018 400046 239558 400102
rect 239614 400046 239682 400102
rect 239738 400046 270278 400102
rect 270334 400046 270402 400102
rect 270458 400046 300998 400102
rect 301054 400046 301122 400102
rect 301178 400046 331718 400102
rect 331774 400046 331842 400102
rect 331898 400046 362438 400102
rect 362494 400046 362562 400102
rect 362618 400046 393158 400102
rect 393214 400046 393282 400102
rect 393338 400046 423878 400102
rect 423934 400046 424002 400102
rect 424058 400046 454598 400102
rect 454654 400046 454722 400102
rect 454778 400046 485318 400102
rect 485374 400046 485442 400102
rect 485498 400046 516038 400102
rect 516094 400046 516162 400102
rect 516218 400046 525250 400102
rect 525306 400046 525374 400102
rect 525430 400046 525498 400102
rect 525554 400046 525622 400102
rect 525678 400046 543250 400102
rect 543306 400046 543374 400102
rect 543430 400046 543498 400102
rect 543554 400046 543622 400102
rect 543678 400046 561250 400102
rect 561306 400046 561374 400102
rect 561430 400046 561498 400102
rect 561554 400046 561622 400102
rect 561678 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 24518 399978
rect 24574 399922 24642 399978
rect 24698 399922 55238 399978
rect 55294 399922 55362 399978
rect 55418 399922 85958 399978
rect 86014 399922 86082 399978
rect 86138 399922 116678 399978
rect 116734 399922 116802 399978
rect 116858 399922 147398 399978
rect 147454 399922 147522 399978
rect 147578 399922 178118 399978
rect 178174 399922 178242 399978
rect 178298 399922 208838 399978
rect 208894 399922 208962 399978
rect 209018 399922 239558 399978
rect 239614 399922 239682 399978
rect 239738 399922 270278 399978
rect 270334 399922 270402 399978
rect 270458 399922 300998 399978
rect 301054 399922 301122 399978
rect 301178 399922 331718 399978
rect 331774 399922 331842 399978
rect 331898 399922 362438 399978
rect 362494 399922 362562 399978
rect 362618 399922 393158 399978
rect 393214 399922 393282 399978
rect 393338 399922 423878 399978
rect 423934 399922 424002 399978
rect 424058 399922 454598 399978
rect 454654 399922 454722 399978
rect 454778 399922 485318 399978
rect 485374 399922 485442 399978
rect 485498 399922 516038 399978
rect 516094 399922 516162 399978
rect 516218 399922 525250 399978
rect 525306 399922 525374 399978
rect 525430 399922 525498 399978
rect 525554 399922 525622 399978
rect 525678 399922 543250 399978
rect 543306 399922 543374 399978
rect 543430 399922 543498 399978
rect 543554 399922 543622 399978
rect 543678 399922 561250 399978
rect 561306 399922 561374 399978
rect 561430 399922 561498 399978
rect 561554 399922 561622 399978
rect 561678 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 39878 388350
rect 39934 388294 40002 388350
rect 40058 388294 70598 388350
rect 70654 388294 70722 388350
rect 70778 388294 101318 388350
rect 101374 388294 101442 388350
rect 101498 388294 132038 388350
rect 132094 388294 132162 388350
rect 132218 388294 162758 388350
rect 162814 388294 162882 388350
rect 162938 388294 193478 388350
rect 193534 388294 193602 388350
rect 193658 388294 224198 388350
rect 224254 388294 224322 388350
rect 224378 388294 254918 388350
rect 254974 388294 255042 388350
rect 255098 388294 285638 388350
rect 285694 388294 285762 388350
rect 285818 388294 316358 388350
rect 316414 388294 316482 388350
rect 316538 388294 347078 388350
rect 347134 388294 347202 388350
rect 347258 388294 377798 388350
rect 377854 388294 377922 388350
rect 377978 388294 408518 388350
rect 408574 388294 408642 388350
rect 408698 388294 439238 388350
rect 439294 388294 439362 388350
rect 439418 388294 469958 388350
rect 470014 388294 470082 388350
rect 470138 388294 500678 388350
rect 500734 388294 500802 388350
rect 500858 388294 528970 388350
rect 529026 388294 529094 388350
rect 529150 388294 529218 388350
rect 529274 388294 529342 388350
rect 529398 388294 546970 388350
rect 547026 388294 547094 388350
rect 547150 388294 547218 388350
rect 547274 388294 547342 388350
rect 547398 388294 564970 388350
rect 565026 388294 565094 388350
rect 565150 388294 565218 388350
rect 565274 388294 565342 388350
rect 565398 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 39878 388226
rect 39934 388170 40002 388226
rect 40058 388170 70598 388226
rect 70654 388170 70722 388226
rect 70778 388170 101318 388226
rect 101374 388170 101442 388226
rect 101498 388170 132038 388226
rect 132094 388170 132162 388226
rect 132218 388170 162758 388226
rect 162814 388170 162882 388226
rect 162938 388170 193478 388226
rect 193534 388170 193602 388226
rect 193658 388170 224198 388226
rect 224254 388170 224322 388226
rect 224378 388170 254918 388226
rect 254974 388170 255042 388226
rect 255098 388170 285638 388226
rect 285694 388170 285762 388226
rect 285818 388170 316358 388226
rect 316414 388170 316482 388226
rect 316538 388170 347078 388226
rect 347134 388170 347202 388226
rect 347258 388170 377798 388226
rect 377854 388170 377922 388226
rect 377978 388170 408518 388226
rect 408574 388170 408642 388226
rect 408698 388170 439238 388226
rect 439294 388170 439362 388226
rect 439418 388170 469958 388226
rect 470014 388170 470082 388226
rect 470138 388170 500678 388226
rect 500734 388170 500802 388226
rect 500858 388170 528970 388226
rect 529026 388170 529094 388226
rect 529150 388170 529218 388226
rect 529274 388170 529342 388226
rect 529398 388170 546970 388226
rect 547026 388170 547094 388226
rect 547150 388170 547218 388226
rect 547274 388170 547342 388226
rect 547398 388170 564970 388226
rect 565026 388170 565094 388226
rect 565150 388170 565218 388226
rect 565274 388170 565342 388226
rect 565398 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 39878 388102
rect 39934 388046 40002 388102
rect 40058 388046 70598 388102
rect 70654 388046 70722 388102
rect 70778 388046 101318 388102
rect 101374 388046 101442 388102
rect 101498 388046 132038 388102
rect 132094 388046 132162 388102
rect 132218 388046 162758 388102
rect 162814 388046 162882 388102
rect 162938 388046 193478 388102
rect 193534 388046 193602 388102
rect 193658 388046 224198 388102
rect 224254 388046 224322 388102
rect 224378 388046 254918 388102
rect 254974 388046 255042 388102
rect 255098 388046 285638 388102
rect 285694 388046 285762 388102
rect 285818 388046 316358 388102
rect 316414 388046 316482 388102
rect 316538 388046 347078 388102
rect 347134 388046 347202 388102
rect 347258 388046 377798 388102
rect 377854 388046 377922 388102
rect 377978 388046 408518 388102
rect 408574 388046 408642 388102
rect 408698 388046 439238 388102
rect 439294 388046 439362 388102
rect 439418 388046 469958 388102
rect 470014 388046 470082 388102
rect 470138 388046 500678 388102
rect 500734 388046 500802 388102
rect 500858 388046 528970 388102
rect 529026 388046 529094 388102
rect 529150 388046 529218 388102
rect 529274 388046 529342 388102
rect 529398 388046 546970 388102
rect 547026 388046 547094 388102
rect 547150 388046 547218 388102
rect 547274 388046 547342 388102
rect 547398 388046 564970 388102
rect 565026 388046 565094 388102
rect 565150 388046 565218 388102
rect 565274 388046 565342 388102
rect 565398 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 39878 387978
rect 39934 387922 40002 387978
rect 40058 387922 70598 387978
rect 70654 387922 70722 387978
rect 70778 387922 101318 387978
rect 101374 387922 101442 387978
rect 101498 387922 132038 387978
rect 132094 387922 132162 387978
rect 132218 387922 162758 387978
rect 162814 387922 162882 387978
rect 162938 387922 193478 387978
rect 193534 387922 193602 387978
rect 193658 387922 224198 387978
rect 224254 387922 224322 387978
rect 224378 387922 254918 387978
rect 254974 387922 255042 387978
rect 255098 387922 285638 387978
rect 285694 387922 285762 387978
rect 285818 387922 316358 387978
rect 316414 387922 316482 387978
rect 316538 387922 347078 387978
rect 347134 387922 347202 387978
rect 347258 387922 377798 387978
rect 377854 387922 377922 387978
rect 377978 387922 408518 387978
rect 408574 387922 408642 387978
rect 408698 387922 439238 387978
rect 439294 387922 439362 387978
rect 439418 387922 469958 387978
rect 470014 387922 470082 387978
rect 470138 387922 500678 387978
rect 500734 387922 500802 387978
rect 500858 387922 528970 387978
rect 529026 387922 529094 387978
rect 529150 387922 529218 387978
rect 529274 387922 529342 387978
rect 529398 387922 546970 387978
rect 547026 387922 547094 387978
rect 547150 387922 547218 387978
rect 547274 387922 547342 387978
rect 547398 387922 564970 387978
rect 565026 387922 565094 387978
rect 565150 387922 565218 387978
rect 565274 387922 565342 387978
rect 565398 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 24518 382350
rect 24574 382294 24642 382350
rect 24698 382294 55238 382350
rect 55294 382294 55362 382350
rect 55418 382294 85958 382350
rect 86014 382294 86082 382350
rect 86138 382294 116678 382350
rect 116734 382294 116802 382350
rect 116858 382294 147398 382350
rect 147454 382294 147522 382350
rect 147578 382294 178118 382350
rect 178174 382294 178242 382350
rect 178298 382294 208838 382350
rect 208894 382294 208962 382350
rect 209018 382294 239558 382350
rect 239614 382294 239682 382350
rect 239738 382294 270278 382350
rect 270334 382294 270402 382350
rect 270458 382294 300998 382350
rect 301054 382294 301122 382350
rect 301178 382294 331718 382350
rect 331774 382294 331842 382350
rect 331898 382294 362438 382350
rect 362494 382294 362562 382350
rect 362618 382294 393158 382350
rect 393214 382294 393282 382350
rect 393338 382294 423878 382350
rect 423934 382294 424002 382350
rect 424058 382294 454598 382350
rect 454654 382294 454722 382350
rect 454778 382294 485318 382350
rect 485374 382294 485442 382350
rect 485498 382294 516038 382350
rect 516094 382294 516162 382350
rect 516218 382294 525250 382350
rect 525306 382294 525374 382350
rect 525430 382294 525498 382350
rect 525554 382294 525622 382350
rect 525678 382294 543250 382350
rect 543306 382294 543374 382350
rect 543430 382294 543498 382350
rect 543554 382294 543622 382350
rect 543678 382294 561250 382350
rect 561306 382294 561374 382350
rect 561430 382294 561498 382350
rect 561554 382294 561622 382350
rect 561678 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 24518 382226
rect 24574 382170 24642 382226
rect 24698 382170 55238 382226
rect 55294 382170 55362 382226
rect 55418 382170 85958 382226
rect 86014 382170 86082 382226
rect 86138 382170 116678 382226
rect 116734 382170 116802 382226
rect 116858 382170 147398 382226
rect 147454 382170 147522 382226
rect 147578 382170 178118 382226
rect 178174 382170 178242 382226
rect 178298 382170 208838 382226
rect 208894 382170 208962 382226
rect 209018 382170 239558 382226
rect 239614 382170 239682 382226
rect 239738 382170 270278 382226
rect 270334 382170 270402 382226
rect 270458 382170 300998 382226
rect 301054 382170 301122 382226
rect 301178 382170 331718 382226
rect 331774 382170 331842 382226
rect 331898 382170 362438 382226
rect 362494 382170 362562 382226
rect 362618 382170 393158 382226
rect 393214 382170 393282 382226
rect 393338 382170 423878 382226
rect 423934 382170 424002 382226
rect 424058 382170 454598 382226
rect 454654 382170 454722 382226
rect 454778 382170 485318 382226
rect 485374 382170 485442 382226
rect 485498 382170 516038 382226
rect 516094 382170 516162 382226
rect 516218 382170 525250 382226
rect 525306 382170 525374 382226
rect 525430 382170 525498 382226
rect 525554 382170 525622 382226
rect 525678 382170 543250 382226
rect 543306 382170 543374 382226
rect 543430 382170 543498 382226
rect 543554 382170 543622 382226
rect 543678 382170 561250 382226
rect 561306 382170 561374 382226
rect 561430 382170 561498 382226
rect 561554 382170 561622 382226
rect 561678 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 24518 382102
rect 24574 382046 24642 382102
rect 24698 382046 55238 382102
rect 55294 382046 55362 382102
rect 55418 382046 85958 382102
rect 86014 382046 86082 382102
rect 86138 382046 116678 382102
rect 116734 382046 116802 382102
rect 116858 382046 147398 382102
rect 147454 382046 147522 382102
rect 147578 382046 178118 382102
rect 178174 382046 178242 382102
rect 178298 382046 208838 382102
rect 208894 382046 208962 382102
rect 209018 382046 239558 382102
rect 239614 382046 239682 382102
rect 239738 382046 270278 382102
rect 270334 382046 270402 382102
rect 270458 382046 300998 382102
rect 301054 382046 301122 382102
rect 301178 382046 331718 382102
rect 331774 382046 331842 382102
rect 331898 382046 362438 382102
rect 362494 382046 362562 382102
rect 362618 382046 393158 382102
rect 393214 382046 393282 382102
rect 393338 382046 423878 382102
rect 423934 382046 424002 382102
rect 424058 382046 454598 382102
rect 454654 382046 454722 382102
rect 454778 382046 485318 382102
rect 485374 382046 485442 382102
rect 485498 382046 516038 382102
rect 516094 382046 516162 382102
rect 516218 382046 525250 382102
rect 525306 382046 525374 382102
rect 525430 382046 525498 382102
rect 525554 382046 525622 382102
rect 525678 382046 543250 382102
rect 543306 382046 543374 382102
rect 543430 382046 543498 382102
rect 543554 382046 543622 382102
rect 543678 382046 561250 382102
rect 561306 382046 561374 382102
rect 561430 382046 561498 382102
rect 561554 382046 561622 382102
rect 561678 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 24518 381978
rect 24574 381922 24642 381978
rect 24698 381922 55238 381978
rect 55294 381922 55362 381978
rect 55418 381922 85958 381978
rect 86014 381922 86082 381978
rect 86138 381922 116678 381978
rect 116734 381922 116802 381978
rect 116858 381922 147398 381978
rect 147454 381922 147522 381978
rect 147578 381922 178118 381978
rect 178174 381922 178242 381978
rect 178298 381922 208838 381978
rect 208894 381922 208962 381978
rect 209018 381922 239558 381978
rect 239614 381922 239682 381978
rect 239738 381922 270278 381978
rect 270334 381922 270402 381978
rect 270458 381922 300998 381978
rect 301054 381922 301122 381978
rect 301178 381922 331718 381978
rect 331774 381922 331842 381978
rect 331898 381922 362438 381978
rect 362494 381922 362562 381978
rect 362618 381922 393158 381978
rect 393214 381922 393282 381978
rect 393338 381922 423878 381978
rect 423934 381922 424002 381978
rect 424058 381922 454598 381978
rect 454654 381922 454722 381978
rect 454778 381922 485318 381978
rect 485374 381922 485442 381978
rect 485498 381922 516038 381978
rect 516094 381922 516162 381978
rect 516218 381922 525250 381978
rect 525306 381922 525374 381978
rect 525430 381922 525498 381978
rect 525554 381922 525622 381978
rect 525678 381922 543250 381978
rect 543306 381922 543374 381978
rect 543430 381922 543498 381978
rect 543554 381922 543622 381978
rect 543678 381922 561250 381978
rect 561306 381922 561374 381978
rect 561430 381922 561498 381978
rect 561554 381922 561622 381978
rect 561678 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 39878 370350
rect 39934 370294 40002 370350
rect 40058 370294 70598 370350
rect 70654 370294 70722 370350
rect 70778 370294 101318 370350
rect 101374 370294 101442 370350
rect 101498 370294 132038 370350
rect 132094 370294 132162 370350
rect 132218 370294 162758 370350
rect 162814 370294 162882 370350
rect 162938 370294 193478 370350
rect 193534 370294 193602 370350
rect 193658 370294 224198 370350
rect 224254 370294 224322 370350
rect 224378 370294 254918 370350
rect 254974 370294 255042 370350
rect 255098 370294 285638 370350
rect 285694 370294 285762 370350
rect 285818 370294 316358 370350
rect 316414 370294 316482 370350
rect 316538 370294 347078 370350
rect 347134 370294 347202 370350
rect 347258 370294 377798 370350
rect 377854 370294 377922 370350
rect 377978 370294 408518 370350
rect 408574 370294 408642 370350
rect 408698 370294 439238 370350
rect 439294 370294 439362 370350
rect 439418 370294 469958 370350
rect 470014 370294 470082 370350
rect 470138 370294 500678 370350
rect 500734 370294 500802 370350
rect 500858 370294 528970 370350
rect 529026 370294 529094 370350
rect 529150 370294 529218 370350
rect 529274 370294 529342 370350
rect 529398 370294 546970 370350
rect 547026 370294 547094 370350
rect 547150 370294 547218 370350
rect 547274 370294 547342 370350
rect 547398 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 39878 370226
rect 39934 370170 40002 370226
rect 40058 370170 70598 370226
rect 70654 370170 70722 370226
rect 70778 370170 101318 370226
rect 101374 370170 101442 370226
rect 101498 370170 132038 370226
rect 132094 370170 132162 370226
rect 132218 370170 162758 370226
rect 162814 370170 162882 370226
rect 162938 370170 193478 370226
rect 193534 370170 193602 370226
rect 193658 370170 224198 370226
rect 224254 370170 224322 370226
rect 224378 370170 254918 370226
rect 254974 370170 255042 370226
rect 255098 370170 285638 370226
rect 285694 370170 285762 370226
rect 285818 370170 316358 370226
rect 316414 370170 316482 370226
rect 316538 370170 347078 370226
rect 347134 370170 347202 370226
rect 347258 370170 377798 370226
rect 377854 370170 377922 370226
rect 377978 370170 408518 370226
rect 408574 370170 408642 370226
rect 408698 370170 439238 370226
rect 439294 370170 439362 370226
rect 439418 370170 469958 370226
rect 470014 370170 470082 370226
rect 470138 370170 500678 370226
rect 500734 370170 500802 370226
rect 500858 370170 528970 370226
rect 529026 370170 529094 370226
rect 529150 370170 529218 370226
rect 529274 370170 529342 370226
rect 529398 370170 546970 370226
rect 547026 370170 547094 370226
rect 547150 370170 547218 370226
rect 547274 370170 547342 370226
rect 547398 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 39878 370102
rect 39934 370046 40002 370102
rect 40058 370046 70598 370102
rect 70654 370046 70722 370102
rect 70778 370046 101318 370102
rect 101374 370046 101442 370102
rect 101498 370046 132038 370102
rect 132094 370046 132162 370102
rect 132218 370046 162758 370102
rect 162814 370046 162882 370102
rect 162938 370046 193478 370102
rect 193534 370046 193602 370102
rect 193658 370046 224198 370102
rect 224254 370046 224322 370102
rect 224378 370046 254918 370102
rect 254974 370046 255042 370102
rect 255098 370046 285638 370102
rect 285694 370046 285762 370102
rect 285818 370046 316358 370102
rect 316414 370046 316482 370102
rect 316538 370046 347078 370102
rect 347134 370046 347202 370102
rect 347258 370046 377798 370102
rect 377854 370046 377922 370102
rect 377978 370046 408518 370102
rect 408574 370046 408642 370102
rect 408698 370046 439238 370102
rect 439294 370046 439362 370102
rect 439418 370046 469958 370102
rect 470014 370046 470082 370102
rect 470138 370046 500678 370102
rect 500734 370046 500802 370102
rect 500858 370046 528970 370102
rect 529026 370046 529094 370102
rect 529150 370046 529218 370102
rect 529274 370046 529342 370102
rect 529398 370046 546970 370102
rect 547026 370046 547094 370102
rect 547150 370046 547218 370102
rect 547274 370046 547342 370102
rect 547398 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 39878 369978
rect 39934 369922 40002 369978
rect 40058 369922 70598 369978
rect 70654 369922 70722 369978
rect 70778 369922 101318 369978
rect 101374 369922 101442 369978
rect 101498 369922 132038 369978
rect 132094 369922 132162 369978
rect 132218 369922 162758 369978
rect 162814 369922 162882 369978
rect 162938 369922 193478 369978
rect 193534 369922 193602 369978
rect 193658 369922 224198 369978
rect 224254 369922 224322 369978
rect 224378 369922 254918 369978
rect 254974 369922 255042 369978
rect 255098 369922 285638 369978
rect 285694 369922 285762 369978
rect 285818 369922 316358 369978
rect 316414 369922 316482 369978
rect 316538 369922 347078 369978
rect 347134 369922 347202 369978
rect 347258 369922 377798 369978
rect 377854 369922 377922 369978
rect 377978 369922 408518 369978
rect 408574 369922 408642 369978
rect 408698 369922 439238 369978
rect 439294 369922 439362 369978
rect 439418 369922 469958 369978
rect 470014 369922 470082 369978
rect 470138 369922 500678 369978
rect 500734 369922 500802 369978
rect 500858 369922 528970 369978
rect 529026 369922 529094 369978
rect 529150 369922 529218 369978
rect 529274 369922 529342 369978
rect 529398 369922 546970 369978
rect 547026 369922 547094 369978
rect 547150 369922 547218 369978
rect 547274 369922 547342 369978
rect 547398 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 24518 364350
rect 24574 364294 24642 364350
rect 24698 364294 55238 364350
rect 55294 364294 55362 364350
rect 55418 364294 85958 364350
rect 86014 364294 86082 364350
rect 86138 364294 116678 364350
rect 116734 364294 116802 364350
rect 116858 364294 147398 364350
rect 147454 364294 147522 364350
rect 147578 364294 178118 364350
rect 178174 364294 178242 364350
rect 178298 364294 208838 364350
rect 208894 364294 208962 364350
rect 209018 364294 239558 364350
rect 239614 364294 239682 364350
rect 239738 364294 270278 364350
rect 270334 364294 270402 364350
rect 270458 364294 300998 364350
rect 301054 364294 301122 364350
rect 301178 364294 331718 364350
rect 331774 364294 331842 364350
rect 331898 364294 362438 364350
rect 362494 364294 362562 364350
rect 362618 364294 393158 364350
rect 393214 364294 393282 364350
rect 393338 364294 423878 364350
rect 423934 364294 424002 364350
rect 424058 364294 454598 364350
rect 454654 364294 454722 364350
rect 454778 364294 485318 364350
rect 485374 364294 485442 364350
rect 485498 364294 516038 364350
rect 516094 364294 516162 364350
rect 516218 364294 525250 364350
rect 525306 364294 525374 364350
rect 525430 364294 525498 364350
rect 525554 364294 525622 364350
rect 525678 364294 543250 364350
rect 543306 364294 543374 364350
rect 543430 364294 543498 364350
rect 543554 364294 543622 364350
rect 543678 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 24518 364226
rect 24574 364170 24642 364226
rect 24698 364170 55238 364226
rect 55294 364170 55362 364226
rect 55418 364170 85958 364226
rect 86014 364170 86082 364226
rect 86138 364170 116678 364226
rect 116734 364170 116802 364226
rect 116858 364170 147398 364226
rect 147454 364170 147522 364226
rect 147578 364170 178118 364226
rect 178174 364170 178242 364226
rect 178298 364170 208838 364226
rect 208894 364170 208962 364226
rect 209018 364170 239558 364226
rect 239614 364170 239682 364226
rect 239738 364170 270278 364226
rect 270334 364170 270402 364226
rect 270458 364170 300998 364226
rect 301054 364170 301122 364226
rect 301178 364170 331718 364226
rect 331774 364170 331842 364226
rect 331898 364170 362438 364226
rect 362494 364170 362562 364226
rect 362618 364170 393158 364226
rect 393214 364170 393282 364226
rect 393338 364170 423878 364226
rect 423934 364170 424002 364226
rect 424058 364170 454598 364226
rect 454654 364170 454722 364226
rect 454778 364170 485318 364226
rect 485374 364170 485442 364226
rect 485498 364170 516038 364226
rect 516094 364170 516162 364226
rect 516218 364170 525250 364226
rect 525306 364170 525374 364226
rect 525430 364170 525498 364226
rect 525554 364170 525622 364226
rect 525678 364170 543250 364226
rect 543306 364170 543374 364226
rect 543430 364170 543498 364226
rect 543554 364170 543622 364226
rect 543678 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 24518 364102
rect 24574 364046 24642 364102
rect 24698 364046 55238 364102
rect 55294 364046 55362 364102
rect 55418 364046 85958 364102
rect 86014 364046 86082 364102
rect 86138 364046 116678 364102
rect 116734 364046 116802 364102
rect 116858 364046 147398 364102
rect 147454 364046 147522 364102
rect 147578 364046 178118 364102
rect 178174 364046 178242 364102
rect 178298 364046 208838 364102
rect 208894 364046 208962 364102
rect 209018 364046 239558 364102
rect 239614 364046 239682 364102
rect 239738 364046 270278 364102
rect 270334 364046 270402 364102
rect 270458 364046 300998 364102
rect 301054 364046 301122 364102
rect 301178 364046 331718 364102
rect 331774 364046 331842 364102
rect 331898 364046 362438 364102
rect 362494 364046 362562 364102
rect 362618 364046 393158 364102
rect 393214 364046 393282 364102
rect 393338 364046 423878 364102
rect 423934 364046 424002 364102
rect 424058 364046 454598 364102
rect 454654 364046 454722 364102
rect 454778 364046 485318 364102
rect 485374 364046 485442 364102
rect 485498 364046 516038 364102
rect 516094 364046 516162 364102
rect 516218 364046 525250 364102
rect 525306 364046 525374 364102
rect 525430 364046 525498 364102
rect 525554 364046 525622 364102
rect 525678 364046 543250 364102
rect 543306 364046 543374 364102
rect 543430 364046 543498 364102
rect 543554 364046 543622 364102
rect 543678 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 24518 363978
rect 24574 363922 24642 363978
rect 24698 363922 55238 363978
rect 55294 363922 55362 363978
rect 55418 363922 85958 363978
rect 86014 363922 86082 363978
rect 86138 363922 116678 363978
rect 116734 363922 116802 363978
rect 116858 363922 147398 363978
rect 147454 363922 147522 363978
rect 147578 363922 178118 363978
rect 178174 363922 178242 363978
rect 178298 363922 208838 363978
rect 208894 363922 208962 363978
rect 209018 363922 239558 363978
rect 239614 363922 239682 363978
rect 239738 363922 270278 363978
rect 270334 363922 270402 363978
rect 270458 363922 300998 363978
rect 301054 363922 301122 363978
rect 301178 363922 331718 363978
rect 331774 363922 331842 363978
rect 331898 363922 362438 363978
rect 362494 363922 362562 363978
rect 362618 363922 393158 363978
rect 393214 363922 393282 363978
rect 393338 363922 423878 363978
rect 423934 363922 424002 363978
rect 424058 363922 454598 363978
rect 454654 363922 454722 363978
rect 454778 363922 485318 363978
rect 485374 363922 485442 363978
rect 485498 363922 516038 363978
rect 516094 363922 516162 363978
rect 516218 363922 525250 363978
rect 525306 363922 525374 363978
rect 525430 363922 525498 363978
rect 525554 363922 525622 363978
rect 525678 363922 543250 363978
rect 543306 363922 543374 363978
rect 543430 363922 543498 363978
rect 543554 363922 543622 363978
rect 543678 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 39878 352350
rect 39934 352294 40002 352350
rect 40058 352294 70598 352350
rect 70654 352294 70722 352350
rect 70778 352294 101318 352350
rect 101374 352294 101442 352350
rect 101498 352294 132038 352350
rect 132094 352294 132162 352350
rect 132218 352294 162758 352350
rect 162814 352294 162882 352350
rect 162938 352294 193478 352350
rect 193534 352294 193602 352350
rect 193658 352294 224198 352350
rect 224254 352294 224322 352350
rect 224378 352294 254918 352350
rect 254974 352294 255042 352350
rect 255098 352294 285638 352350
rect 285694 352294 285762 352350
rect 285818 352294 316358 352350
rect 316414 352294 316482 352350
rect 316538 352294 347078 352350
rect 347134 352294 347202 352350
rect 347258 352294 377798 352350
rect 377854 352294 377922 352350
rect 377978 352294 408518 352350
rect 408574 352294 408642 352350
rect 408698 352294 439238 352350
rect 439294 352294 439362 352350
rect 439418 352294 469958 352350
rect 470014 352294 470082 352350
rect 470138 352294 500678 352350
rect 500734 352294 500802 352350
rect 500858 352294 528970 352350
rect 529026 352294 529094 352350
rect 529150 352294 529218 352350
rect 529274 352294 529342 352350
rect 529398 352294 546970 352350
rect 547026 352294 547094 352350
rect 547150 352294 547218 352350
rect 547274 352294 547342 352350
rect 547398 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 39878 352226
rect 39934 352170 40002 352226
rect 40058 352170 70598 352226
rect 70654 352170 70722 352226
rect 70778 352170 101318 352226
rect 101374 352170 101442 352226
rect 101498 352170 132038 352226
rect 132094 352170 132162 352226
rect 132218 352170 162758 352226
rect 162814 352170 162882 352226
rect 162938 352170 193478 352226
rect 193534 352170 193602 352226
rect 193658 352170 224198 352226
rect 224254 352170 224322 352226
rect 224378 352170 254918 352226
rect 254974 352170 255042 352226
rect 255098 352170 285638 352226
rect 285694 352170 285762 352226
rect 285818 352170 316358 352226
rect 316414 352170 316482 352226
rect 316538 352170 347078 352226
rect 347134 352170 347202 352226
rect 347258 352170 377798 352226
rect 377854 352170 377922 352226
rect 377978 352170 408518 352226
rect 408574 352170 408642 352226
rect 408698 352170 439238 352226
rect 439294 352170 439362 352226
rect 439418 352170 469958 352226
rect 470014 352170 470082 352226
rect 470138 352170 500678 352226
rect 500734 352170 500802 352226
rect 500858 352170 528970 352226
rect 529026 352170 529094 352226
rect 529150 352170 529218 352226
rect 529274 352170 529342 352226
rect 529398 352170 546970 352226
rect 547026 352170 547094 352226
rect 547150 352170 547218 352226
rect 547274 352170 547342 352226
rect 547398 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 39878 352102
rect 39934 352046 40002 352102
rect 40058 352046 70598 352102
rect 70654 352046 70722 352102
rect 70778 352046 101318 352102
rect 101374 352046 101442 352102
rect 101498 352046 132038 352102
rect 132094 352046 132162 352102
rect 132218 352046 162758 352102
rect 162814 352046 162882 352102
rect 162938 352046 193478 352102
rect 193534 352046 193602 352102
rect 193658 352046 224198 352102
rect 224254 352046 224322 352102
rect 224378 352046 254918 352102
rect 254974 352046 255042 352102
rect 255098 352046 285638 352102
rect 285694 352046 285762 352102
rect 285818 352046 316358 352102
rect 316414 352046 316482 352102
rect 316538 352046 347078 352102
rect 347134 352046 347202 352102
rect 347258 352046 377798 352102
rect 377854 352046 377922 352102
rect 377978 352046 408518 352102
rect 408574 352046 408642 352102
rect 408698 352046 439238 352102
rect 439294 352046 439362 352102
rect 439418 352046 469958 352102
rect 470014 352046 470082 352102
rect 470138 352046 500678 352102
rect 500734 352046 500802 352102
rect 500858 352046 528970 352102
rect 529026 352046 529094 352102
rect 529150 352046 529218 352102
rect 529274 352046 529342 352102
rect 529398 352046 546970 352102
rect 547026 352046 547094 352102
rect 547150 352046 547218 352102
rect 547274 352046 547342 352102
rect 547398 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 39878 351978
rect 39934 351922 40002 351978
rect 40058 351922 70598 351978
rect 70654 351922 70722 351978
rect 70778 351922 101318 351978
rect 101374 351922 101442 351978
rect 101498 351922 132038 351978
rect 132094 351922 132162 351978
rect 132218 351922 162758 351978
rect 162814 351922 162882 351978
rect 162938 351922 193478 351978
rect 193534 351922 193602 351978
rect 193658 351922 224198 351978
rect 224254 351922 224322 351978
rect 224378 351922 254918 351978
rect 254974 351922 255042 351978
rect 255098 351922 285638 351978
rect 285694 351922 285762 351978
rect 285818 351922 316358 351978
rect 316414 351922 316482 351978
rect 316538 351922 347078 351978
rect 347134 351922 347202 351978
rect 347258 351922 377798 351978
rect 377854 351922 377922 351978
rect 377978 351922 408518 351978
rect 408574 351922 408642 351978
rect 408698 351922 439238 351978
rect 439294 351922 439362 351978
rect 439418 351922 469958 351978
rect 470014 351922 470082 351978
rect 470138 351922 500678 351978
rect 500734 351922 500802 351978
rect 500858 351922 528970 351978
rect 529026 351922 529094 351978
rect 529150 351922 529218 351978
rect 529274 351922 529342 351978
rect 529398 351922 546970 351978
rect 547026 351922 547094 351978
rect 547150 351922 547218 351978
rect 547274 351922 547342 351978
rect 547398 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 24518 346350
rect 24574 346294 24642 346350
rect 24698 346294 55238 346350
rect 55294 346294 55362 346350
rect 55418 346294 85958 346350
rect 86014 346294 86082 346350
rect 86138 346294 116678 346350
rect 116734 346294 116802 346350
rect 116858 346294 147398 346350
rect 147454 346294 147522 346350
rect 147578 346294 178118 346350
rect 178174 346294 178242 346350
rect 178298 346294 208838 346350
rect 208894 346294 208962 346350
rect 209018 346294 239558 346350
rect 239614 346294 239682 346350
rect 239738 346294 270278 346350
rect 270334 346294 270402 346350
rect 270458 346294 300998 346350
rect 301054 346294 301122 346350
rect 301178 346294 331718 346350
rect 331774 346294 331842 346350
rect 331898 346294 362438 346350
rect 362494 346294 362562 346350
rect 362618 346294 393158 346350
rect 393214 346294 393282 346350
rect 393338 346294 423878 346350
rect 423934 346294 424002 346350
rect 424058 346294 454598 346350
rect 454654 346294 454722 346350
rect 454778 346294 485318 346350
rect 485374 346294 485442 346350
rect 485498 346294 516038 346350
rect 516094 346294 516162 346350
rect 516218 346294 525250 346350
rect 525306 346294 525374 346350
rect 525430 346294 525498 346350
rect 525554 346294 525622 346350
rect 525678 346294 543250 346350
rect 543306 346294 543374 346350
rect 543430 346294 543498 346350
rect 543554 346294 543622 346350
rect 543678 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 24518 346226
rect 24574 346170 24642 346226
rect 24698 346170 55238 346226
rect 55294 346170 55362 346226
rect 55418 346170 85958 346226
rect 86014 346170 86082 346226
rect 86138 346170 116678 346226
rect 116734 346170 116802 346226
rect 116858 346170 147398 346226
rect 147454 346170 147522 346226
rect 147578 346170 178118 346226
rect 178174 346170 178242 346226
rect 178298 346170 208838 346226
rect 208894 346170 208962 346226
rect 209018 346170 239558 346226
rect 239614 346170 239682 346226
rect 239738 346170 270278 346226
rect 270334 346170 270402 346226
rect 270458 346170 300998 346226
rect 301054 346170 301122 346226
rect 301178 346170 331718 346226
rect 331774 346170 331842 346226
rect 331898 346170 362438 346226
rect 362494 346170 362562 346226
rect 362618 346170 393158 346226
rect 393214 346170 393282 346226
rect 393338 346170 423878 346226
rect 423934 346170 424002 346226
rect 424058 346170 454598 346226
rect 454654 346170 454722 346226
rect 454778 346170 485318 346226
rect 485374 346170 485442 346226
rect 485498 346170 516038 346226
rect 516094 346170 516162 346226
rect 516218 346170 525250 346226
rect 525306 346170 525374 346226
rect 525430 346170 525498 346226
rect 525554 346170 525622 346226
rect 525678 346170 543250 346226
rect 543306 346170 543374 346226
rect 543430 346170 543498 346226
rect 543554 346170 543622 346226
rect 543678 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 24518 346102
rect 24574 346046 24642 346102
rect 24698 346046 55238 346102
rect 55294 346046 55362 346102
rect 55418 346046 85958 346102
rect 86014 346046 86082 346102
rect 86138 346046 116678 346102
rect 116734 346046 116802 346102
rect 116858 346046 147398 346102
rect 147454 346046 147522 346102
rect 147578 346046 178118 346102
rect 178174 346046 178242 346102
rect 178298 346046 208838 346102
rect 208894 346046 208962 346102
rect 209018 346046 239558 346102
rect 239614 346046 239682 346102
rect 239738 346046 270278 346102
rect 270334 346046 270402 346102
rect 270458 346046 300998 346102
rect 301054 346046 301122 346102
rect 301178 346046 331718 346102
rect 331774 346046 331842 346102
rect 331898 346046 362438 346102
rect 362494 346046 362562 346102
rect 362618 346046 393158 346102
rect 393214 346046 393282 346102
rect 393338 346046 423878 346102
rect 423934 346046 424002 346102
rect 424058 346046 454598 346102
rect 454654 346046 454722 346102
rect 454778 346046 485318 346102
rect 485374 346046 485442 346102
rect 485498 346046 516038 346102
rect 516094 346046 516162 346102
rect 516218 346046 525250 346102
rect 525306 346046 525374 346102
rect 525430 346046 525498 346102
rect 525554 346046 525622 346102
rect 525678 346046 543250 346102
rect 543306 346046 543374 346102
rect 543430 346046 543498 346102
rect 543554 346046 543622 346102
rect 543678 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 24518 345978
rect 24574 345922 24642 345978
rect 24698 345922 55238 345978
rect 55294 345922 55362 345978
rect 55418 345922 85958 345978
rect 86014 345922 86082 345978
rect 86138 345922 116678 345978
rect 116734 345922 116802 345978
rect 116858 345922 147398 345978
rect 147454 345922 147522 345978
rect 147578 345922 178118 345978
rect 178174 345922 178242 345978
rect 178298 345922 208838 345978
rect 208894 345922 208962 345978
rect 209018 345922 239558 345978
rect 239614 345922 239682 345978
rect 239738 345922 270278 345978
rect 270334 345922 270402 345978
rect 270458 345922 300998 345978
rect 301054 345922 301122 345978
rect 301178 345922 331718 345978
rect 331774 345922 331842 345978
rect 331898 345922 362438 345978
rect 362494 345922 362562 345978
rect 362618 345922 393158 345978
rect 393214 345922 393282 345978
rect 393338 345922 423878 345978
rect 423934 345922 424002 345978
rect 424058 345922 454598 345978
rect 454654 345922 454722 345978
rect 454778 345922 485318 345978
rect 485374 345922 485442 345978
rect 485498 345922 516038 345978
rect 516094 345922 516162 345978
rect 516218 345922 525250 345978
rect 525306 345922 525374 345978
rect 525430 345922 525498 345978
rect 525554 345922 525622 345978
rect 525678 345922 543250 345978
rect 543306 345922 543374 345978
rect 543430 345922 543498 345978
rect 543554 345922 543622 345978
rect 543678 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 39878 334350
rect 39934 334294 40002 334350
rect 40058 334294 70598 334350
rect 70654 334294 70722 334350
rect 70778 334294 101318 334350
rect 101374 334294 101442 334350
rect 101498 334294 132038 334350
rect 132094 334294 132162 334350
rect 132218 334294 162758 334350
rect 162814 334294 162882 334350
rect 162938 334294 193478 334350
rect 193534 334294 193602 334350
rect 193658 334294 224198 334350
rect 224254 334294 224322 334350
rect 224378 334294 254918 334350
rect 254974 334294 255042 334350
rect 255098 334294 285638 334350
rect 285694 334294 285762 334350
rect 285818 334294 316358 334350
rect 316414 334294 316482 334350
rect 316538 334294 347078 334350
rect 347134 334294 347202 334350
rect 347258 334294 377798 334350
rect 377854 334294 377922 334350
rect 377978 334294 408518 334350
rect 408574 334294 408642 334350
rect 408698 334294 439238 334350
rect 439294 334294 439362 334350
rect 439418 334294 469958 334350
rect 470014 334294 470082 334350
rect 470138 334294 500678 334350
rect 500734 334294 500802 334350
rect 500858 334294 528970 334350
rect 529026 334294 529094 334350
rect 529150 334294 529218 334350
rect 529274 334294 529342 334350
rect 529398 334294 546970 334350
rect 547026 334294 547094 334350
rect 547150 334294 547218 334350
rect 547274 334294 547342 334350
rect 547398 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 39878 334226
rect 39934 334170 40002 334226
rect 40058 334170 70598 334226
rect 70654 334170 70722 334226
rect 70778 334170 101318 334226
rect 101374 334170 101442 334226
rect 101498 334170 132038 334226
rect 132094 334170 132162 334226
rect 132218 334170 162758 334226
rect 162814 334170 162882 334226
rect 162938 334170 193478 334226
rect 193534 334170 193602 334226
rect 193658 334170 224198 334226
rect 224254 334170 224322 334226
rect 224378 334170 254918 334226
rect 254974 334170 255042 334226
rect 255098 334170 285638 334226
rect 285694 334170 285762 334226
rect 285818 334170 316358 334226
rect 316414 334170 316482 334226
rect 316538 334170 347078 334226
rect 347134 334170 347202 334226
rect 347258 334170 377798 334226
rect 377854 334170 377922 334226
rect 377978 334170 408518 334226
rect 408574 334170 408642 334226
rect 408698 334170 439238 334226
rect 439294 334170 439362 334226
rect 439418 334170 469958 334226
rect 470014 334170 470082 334226
rect 470138 334170 500678 334226
rect 500734 334170 500802 334226
rect 500858 334170 528970 334226
rect 529026 334170 529094 334226
rect 529150 334170 529218 334226
rect 529274 334170 529342 334226
rect 529398 334170 546970 334226
rect 547026 334170 547094 334226
rect 547150 334170 547218 334226
rect 547274 334170 547342 334226
rect 547398 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 39878 334102
rect 39934 334046 40002 334102
rect 40058 334046 70598 334102
rect 70654 334046 70722 334102
rect 70778 334046 101318 334102
rect 101374 334046 101442 334102
rect 101498 334046 132038 334102
rect 132094 334046 132162 334102
rect 132218 334046 162758 334102
rect 162814 334046 162882 334102
rect 162938 334046 193478 334102
rect 193534 334046 193602 334102
rect 193658 334046 224198 334102
rect 224254 334046 224322 334102
rect 224378 334046 254918 334102
rect 254974 334046 255042 334102
rect 255098 334046 285638 334102
rect 285694 334046 285762 334102
rect 285818 334046 316358 334102
rect 316414 334046 316482 334102
rect 316538 334046 347078 334102
rect 347134 334046 347202 334102
rect 347258 334046 377798 334102
rect 377854 334046 377922 334102
rect 377978 334046 408518 334102
rect 408574 334046 408642 334102
rect 408698 334046 439238 334102
rect 439294 334046 439362 334102
rect 439418 334046 469958 334102
rect 470014 334046 470082 334102
rect 470138 334046 500678 334102
rect 500734 334046 500802 334102
rect 500858 334046 528970 334102
rect 529026 334046 529094 334102
rect 529150 334046 529218 334102
rect 529274 334046 529342 334102
rect 529398 334046 546970 334102
rect 547026 334046 547094 334102
rect 547150 334046 547218 334102
rect 547274 334046 547342 334102
rect 547398 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 39878 333978
rect 39934 333922 40002 333978
rect 40058 333922 70598 333978
rect 70654 333922 70722 333978
rect 70778 333922 101318 333978
rect 101374 333922 101442 333978
rect 101498 333922 132038 333978
rect 132094 333922 132162 333978
rect 132218 333922 162758 333978
rect 162814 333922 162882 333978
rect 162938 333922 193478 333978
rect 193534 333922 193602 333978
rect 193658 333922 224198 333978
rect 224254 333922 224322 333978
rect 224378 333922 254918 333978
rect 254974 333922 255042 333978
rect 255098 333922 285638 333978
rect 285694 333922 285762 333978
rect 285818 333922 316358 333978
rect 316414 333922 316482 333978
rect 316538 333922 347078 333978
rect 347134 333922 347202 333978
rect 347258 333922 377798 333978
rect 377854 333922 377922 333978
rect 377978 333922 408518 333978
rect 408574 333922 408642 333978
rect 408698 333922 439238 333978
rect 439294 333922 439362 333978
rect 439418 333922 469958 333978
rect 470014 333922 470082 333978
rect 470138 333922 500678 333978
rect 500734 333922 500802 333978
rect 500858 333922 528970 333978
rect 529026 333922 529094 333978
rect 529150 333922 529218 333978
rect 529274 333922 529342 333978
rect 529398 333922 546970 333978
rect 547026 333922 547094 333978
rect 547150 333922 547218 333978
rect 547274 333922 547342 333978
rect 547398 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 24518 328350
rect 24574 328294 24642 328350
rect 24698 328294 55238 328350
rect 55294 328294 55362 328350
rect 55418 328294 85958 328350
rect 86014 328294 86082 328350
rect 86138 328294 116678 328350
rect 116734 328294 116802 328350
rect 116858 328294 147398 328350
rect 147454 328294 147522 328350
rect 147578 328294 178118 328350
rect 178174 328294 178242 328350
rect 178298 328294 208838 328350
rect 208894 328294 208962 328350
rect 209018 328294 239558 328350
rect 239614 328294 239682 328350
rect 239738 328294 270278 328350
rect 270334 328294 270402 328350
rect 270458 328294 300998 328350
rect 301054 328294 301122 328350
rect 301178 328294 331718 328350
rect 331774 328294 331842 328350
rect 331898 328294 362438 328350
rect 362494 328294 362562 328350
rect 362618 328294 393158 328350
rect 393214 328294 393282 328350
rect 393338 328294 423878 328350
rect 423934 328294 424002 328350
rect 424058 328294 454598 328350
rect 454654 328294 454722 328350
rect 454778 328294 485318 328350
rect 485374 328294 485442 328350
rect 485498 328294 516038 328350
rect 516094 328294 516162 328350
rect 516218 328294 525250 328350
rect 525306 328294 525374 328350
rect 525430 328294 525498 328350
rect 525554 328294 525622 328350
rect 525678 328294 543250 328350
rect 543306 328294 543374 328350
rect 543430 328294 543498 328350
rect 543554 328294 543622 328350
rect 543678 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 24518 328226
rect 24574 328170 24642 328226
rect 24698 328170 55238 328226
rect 55294 328170 55362 328226
rect 55418 328170 85958 328226
rect 86014 328170 86082 328226
rect 86138 328170 116678 328226
rect 116734 328170 116802 328226
rect 116858 328170 147398 328226
rect 147454 328170 147522 328226
rect 147578 328170 178118 328226
rect 178174 328170 178242 328226
rect 178298 328170 208838 328226
rect 208894 328170 208962 328226
rect 209018 328170 239558 328226
rect 239614 328170 239682 328226
rect 239738 328170 270278 328226
rect 270334 328170 270402 328226
rect 270458 328170 300998 328226
rect 301054 328170 301122 328226
rect 301178 328170 331718 328226
rect 331774 328170 331842 328226
rect 331898 328170 362438 328226
rect 362494 328170 362562 328226
rect 362618 328170 393158 328226
rect 393214 328170 393282 328226
rect 393338 328170 423878 328226
rect 423934 328170 424002 328226
rect 424058 328170 454598 328226
rect 454654 328170 454722 328226
rect 454778 328170 485318 328226
rect 485374 328170 485442 328226
rect 485498 328170 516038 328226
rect 516094 328170 516162 328226
rect 516218 328170 525250 328226
rect 525306 328170 525374 328226
rect 525430 328170 525498 328226
rect 525554 328170 525622 328226
rect 525678 328170 543250 328226
rect 543306 328170 543374 328226
rect 543430 328170 543498 328226
rect 543554 328170 543622 328226
rect 543678 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 24518 328102
rect 24574 328046 24642 328102
rect 24698 328046 55238 328102
rect 55294 328046 55362 328102
rect 55418 328046 85958 328102
rect 86014 328046 86082 328102
rect 86138 328046 116678 328102
rect 116734 328046 116802 328102
rect 116858 328046 147398 328102
rect 147454 328046 147522 328102
rect 147578 328046 178118 328102
rect 178174 328046 178242 328102
rect 178298 328046 208838 328102
rect 208894 328046 208962 328102
rect 209018 328046 239558 328102
rect 239614 328046 239682 328102
rect 239738 328046 270278 328102
rect 270334 328046 270402 328102
rect 270458 328046 300998 328102
rect 301054 328046 301122 328102
rect 301178 328046 331718 328102
rect 331774 328046 331842 328102
rect 331898 328046 362438 328102
rect 362494 328046 362562 328102
rect 362618 328046 393158 328102
rect 393214 328046 393282 328102
rect 393338 328046 423878 328102
rect 423934 328046 424002 328102
rect 424058 328046 454598 328102
rect 454654 328046 454722 328102
rect 454778 328046 485318 328102
rect 485374 328046 485442 328102
rect 485498 328046 516038 328102
rect 516094 328046 516162 328102
rect 516218 328046 525250 328102
rect 525306 328046 525374 328102
rect 525430 328046 525498 328102
rect 525554 328046 525622 328102
rect 525678 328046 543250 328102
rect 543306 328046 543374 328102
rect 543430 328046 543498 328102
rect 543554 328046 543622 328102
rect 543678 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 24518 327978
rect 24574 327922 24642 327978
rect 24698 327922 55238 327978
rect 55294 327922 55362 327978
rect 55418 327922 85958 327978
rect 86014 327922 86082 327978
rect 86138 327922 116678 327978
rect 116734 327922 116802 327978
rect 116858 327922 147398 327978
rect 147454 327922 147522 327978
rect 147578 327922 178118 327978
rect 178174 327922 178242 327978
rect 178298 327922 208838 327978
rect 208894 327922 208962 327978
rect 209018 327922 239558 327978
rect 239614 327922 239682 327978
rect 239738 327922 270278 327978
rect 270334 327922 270402 327978
rect 270458 327922 300998 327978
rect 301054 327922 301122 327978
rect 301178 327922 331718 327978
rect 331774 327922 331842 327978
rect 331898 327922 362438 327978
rect 362494 327922 362562 327978
rect 362618 327922 393158 327978
rect 393214 327922 393282 327978
rect 393338 327922 423878 327978
rect 423934 327922 424002 327978
rect 424058 327922 454598 327978
rect 454654 327922 454722 327978
rect 454778 327922 485318 327978
rect 485374 327922 485442 327978
rect 485498 327922 516038 327978
rect 516094 327922 516162 327978
rect 516218 327922 525250 327978
rect 525306 327922 525374 327978
rect 525430 327922 525498 327978
rect 525554 327922 525622 327978
rect 525678 327922 543250 327978
rect 543306 327922 543374 327978
rect 543430 327922 543498 327978
rect 543554 327922 543622 327978
rect 543678 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 39878 316350
rect 39934 316294 40002 316350
rect 40058 316294 70598 316350
rect 70654 316294 70722 316350
rect 70778 316294 101318 316350
rect 101374 316294 101442 316350
rect 101498 316294 132038 316350
rect 132094 316294 132162 316350
rect 132218 316294 162758 316350
rect 162814 316294 162882 316350
rect 162938 316294 193478 316350
rect 193534 316294 193602 316350
rect 193658 316294 224198 316350
rect 224254 316294 224322 316350
rect 224378 316294 254918 316350
rect 254974 316294 255042 316350
rect 255098 316294 285638 316350
rect 285694 316294 285762 316350
rect 285818 316294 316358 316350
rect 316414 316294 316482 316350
rect 316538 316294 347078 316350
rect 347134 316294 347202 316350
rect 347258 316294 377798 316350
rect 377854 316294 377922 316350
rect 377978 316294 408518 316350
rect 408574 316294 408642 316350
rect 408698 316294 439238 316350
rect 439294 316294 439362 316350
rect 439418 316294 469958 316350
rect 470014 316294 470082 316350
rect 470138 316294 500678 316350
rect 500734 316294 500802 316350
rect 500858 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 39878 316226
rect 39934 316170 40002 316226
rect 40058 316170 70598 316226
rect 70654 316170 70722 316226
rect 70778 316170 101318 316226
rect 101374 316170 101442 316226
rect 101498 316170 132038 316226
rect 132094 316170 132162 316226
rect 132218 316170 162758 316226
rect 162814 316170 162882 316226
rect 162938 316170 193478 316226
rect 193534 316170 193602 316226
rect 193658 316170 224198 316226
rect 224254 316170 224322 316226
rect 224378 316170 254918 316226
rect 254974 316170 255042 316226
rect 255098 316170 285638 316226
rect 285694 316170 285762 316226
rect 285818 316170 316358 316226
rect 316414 316170 316482 316226
rect 316538 316170 347078 316226
rect 347134 316170 347202 316226
rect 347258 316170 377798 316226
rect 377854 316170 377922 316226
rect 377978 316170 408518 316226
rect 408574 316170 408642 316226
rect 408698 316170 439238 316226
rect 439294 316170 439362 316226
rect 439418 316170 469958 316226
rect 470014 316170 470082 316226
rect 470138 316170 500678 316226
rect 500734 316170 500802 316226
rect 500858 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 39878 316102
rect 39934 316046 40002 316102
rect 40058 316046 70598 316102
rect 70654 316046 70722 316102
rect 70778 316046 101318 316102
rect 101374 316046 101442 316102
rect 101498 316046 132038 316102
rect 132094 316046 132162 316102
rect 132218 316046 162758 316102
rect 162814 316046 162882 316102
rect 162938 316046 193478 316102
rect 193534 316046 193602 316102
rect 193658 316046 224198 316102
rect 224254 316046 224322 316102
rect 224378 316046 254918 316102
rect 254974 316046 255042 316102
rect 255098 316046 285638 316102
rect 285694 316046 285762 316102
rect 285818 316046 316358 316102
rect 316414 316046 316482 316102
rect 316538 316046 347078 316102
rect 347134 316046 347202 316102
rect 347258 316046 377798 316102
rect 377854 316046 377922 316102
rect 377978 316046 408518 316102
rect 408574 316046 408642 316102
rect 408698 316046 439238 316102
rect 439294 316046 439362 316102
rect 439418 316046 469958 316102
rect 470014 316046 470082 316102
rect 470138 316046 500678 316102
rect 500734 316046 500802 316102
rect 500858 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 39878 315978
rect 39934 315922 40002 315978
rect 40058 315922 70598 315978
rect 70654 315922 70722 315978
rect 70778 315922 101318 315978
rect 101374 315922 101442 315978
rect 101498 315922 132038 315978
rect 132094 315922 132162 315978
rect 132218 315922 162758 315978
rect 162814 315922 162882 315978
rect 162938 315922 193478 315978
rect 193534 315922 193602 315978
rect 193658 315922 224198 315978
rect 224254 315922 224322 315978
rect 224378 315922 254918 315978
rect 254974 315922 255042 315978
rect 255098 315922 285638 315978
rect 285694 315922 285762 315978
rect 285818 315922 316358 315978
rect 316414 315922 316482 315978
rect 316538 315922 347078 315978
rect 347134 315922 347202 315978
rect 347258 315922 377798 315978
rect 377854 315922 377922 315978
rect 377978 315922 408518 315978
rect 408574 315922 408642 315978
rect 408698 315922 439238 315978
rect 439294 315922 439362 315978
rect 439418 315922 469958 315978
rect 470014 315922 470082 315978
rect 470138 315922 500678 315978
rect 500734 315922 500802 315978
rect 500858 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 24518 310350
rect 24574 310294 24642 310350
rect 24698 310294 55238 310350
rect 55294 310294 55362 310350
rect 55418 310294 85958 310350
rect 86014 310294 86082 310350
rect 86138 310294 116678 310350
rect 116734 310294 116802 310350
rect 116858 310294 147398 310350
rect 147454 310294 147522 310350
rect 147578 310294 178118 310350
rect 178174 310294 178242 310350
rect 178298 310294 208838 310350
rect 208894 310294 208962 310350
rect 209018 310294 239558 310350
rect 239614 310294 239682 310350
rect 239738 310294 270278 310350
rect 270334 310294 270402 310350
rect 270458 310294 300998 310350
rect 301054 310294 301122 310350
rect 301178 310294 331718 310350
rect 331774 310294 331842 310350
rect 331898 310294 362438 310350
rect 362494 310294 362562 310350
rect 362618 310294 393158 310350
rect 393214 310294 393282 310350
rect 393338 310294 423878 310350
rect 423934 310294 424002 310350
rect 424058 310294 454598 310350
rect 454654 310294 454722 310350
rect 454778 310294 485318 310350
rect 485374 310294 485442 310350
rect 485498 310294 516038 310350
rect 516094 310294 516162 310350
rect 516218 310294 525250 310350
rect 525306 310294 525374 310350
rect 525430 310294 525498 310350
rect 525554 310294 525622 310350
rect 525678 310294 543250 310350
rect 543306 310294 543374 310350
rect 543430 310294 543498 310350
rect 543554 310294 543622 310350
rect 543678 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 24518 310226
rect 24574 310170 24642 310226
rect 24698 310170 55238 310226
rect 55294 310170 55362 310226
rect 55418 310170 85958 310226
rect 86014 310170 86082 310226
rect 86138 310170 116678 310226
rect 116734 310170 116802 310226
rect 116858 310170 147398 310226
rect 147454 310170 147522 310226
rect 147578 310170 178118 310226
rect 178174 310170 178242 310226
rect 178298 310170 208838 310226
rect 208894 310170 208962 310226
rect 209018 310170 239558 310226
rect 239614 310170 239682 310226
rect 239738 310170 270278 310226
rect 270334 310170 270402 310226
rect 270458 310170 300998 310226
rect 301054 310170 301122 310226
rect 301178 310170 331718 310226
rect 331774 310170 331842 310226
rect 331898 310170 362438 310226
rect 362494 310170 362562 310226
rect 362618 310170 393158 310226
rect 393214 310170 393282 310226
rect 393338 310170 423878 310226
rect 423934 310170 424002 310226
rect 424058 310170 454598 310226
rect 454654 310170 454722 310226
rect 454778 310170 485318 310226
rect 485374 310170 485442 310226
rect 485498 310170 516038 310226
rect 516094 310170 516162 310226
rect 516218 310170 525250 310226
rect 525306 310170 525374 310226
rect 525430 310170 525498 310226
rect 525554 310170 525622 310226
rect 525678 310170 543250 310226
rect 543306 310170 543374 310226
rect 543430 310170 543498 310226
rect 543554 310170 543622 310226
rect 543678 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 24518 310102
rect 24574 310046 24642 310102
rect 24698 310046 55238 310102
rect 55294 310046 55362 310102
rect 55418 310046 85958 310102
rect 86014 310046 86082 310102
rect 86138 310046 116678 310102
rect 116734 310046 116802 310102
rect 116858 310046 147398 310102
rect 147454 310046 147522 310102
rect 147578 310046 178118 310102
rect 178174 310046 178242 310102
rect 178298 310046 208838 310102
rect 208894 310046 208962 310102
rect 209018 310046 239558 310102
rect 239614 310046 239682 310102
rect 239738 310046 270278 310102
rect 270334 310046 270402 310102
rect 270458 310046 300998 310102
rect 301054 310046 301122 310102
rect 301178 310046 331718 310102
rect 331774 310046 331842 310102
rect 331898 310046 362438 310102
rect 362494 310046 362562 310102
rect 362618 310046 393158 310102
rect 393214 310046 393282 310102
rect 393338 310046 423878 310102
rect 423934 310046 424002 310102
rect 424058 310046 454598 310102
rect 454654 310046 454722 310102
rect 454778 310046 485318 310102
rect 485374 310046 485442 310102
rect 485498 310046 516038 310102
rect 516094 310046 516162 310102
rect 516218 310046 525250 310102
rect 525306 310046 525374 310102
rect 525430 310046 525498 310102
rect 525554 310046 525622 310102
rect 525678 310046 543250 310102
rect 543306 310046 543374 310102
rect 543430 310046 543498 310102
rect 543554 310046 543622 310102
rect 543678 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 24518 309978
rect 24574 309922 24642 309978
rect 24698 309922 55238 309978
rect 55294 309922 55362 309978
rect 55418 309922 85958 309978
rect 86014 309922 86082 309978
rect 86138 309922 116678 309978
rect 116734 309922 116802 309978
rect 116858 309922 147398 309978
rect 147454 309922 147522 309978
rect 147578 309922 178118 309978
rect 178174 309922 178242 309978
rect 178298 309922 208838 309978
rect 208894 309922 208962 309978
rect 209018 309922 239558 309978
rect 239614 309922 239682 309978
rect 239738 309922 270278 309978
rect 270334 309922 270402 309978
rect 270458 309922 300998 309978
rect 301054 309922 301122 309978
rect 301178 309922 331718 309978
rect 331774 309922 331842 309978
rect 331898 309922 362438 309978
rect 362494 309922 362562 309978
rect 362618 309922 393158 309978
rect 393214 309922 393282 309978
rect 393338 309922 423878 309978
rect 423934 309922 424002 309978
rect 424058 309922 454598 309978
rect 454654 309922 454722 309978
rect 454778 309922 485318 309978
rect 485374 309922 485442 309978
rect 485498 309922 516038 309978
rect 516094 309922 516162 309978
rect 516218 309922 525250 309978
rect 525306 309922 525374 309978
rect 525430 309922 525498 309978
rect 525554 309922 525622 309978
rect 525678 309922 543250 309978
rect 543306 309922 543374 309978
rect 543430 309922 543498 309978
rect 543554 309922 543622 309978
rect 543678 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 39878 298350
rect 39934 298294 40002 298350
rect 40058 298294 70598 298350
rect 70654 298294 70722 298350
rect 70778 298294 101318 298350
rect 101374 298294 101442 298350
rect 101498 298294 132038 298350
rect 132094 298294 132162 298350
rect 132218 298294 162758 298350
rect 162814 298294 162882 298350
rect 162938 298294 193478 298350
rect 193534 298294 193602 298350
rect 193658 298294 224198 298350
rect 224254 298294 224322 298350
rect 224378 298294 254918 298350
rect 254974 298294 255042 298350
rect 255098 298294 285638 298350
rect 285694 298294 285762 298350
rect 285818 298294 316358 298350
rect 316414 298294 316482 298350
rect 316538 298294 347078 298350
rect 347134 298294 347202 298350
rect 347258 298294 377798 298350
rect 377854 298294 377922 298350
rect 377978 298294 408518 298350
rect 408574 298294 408642 298350
rect 408698 298294 439238 298350
rect 439294 298294 439362 298350
rect 439418 298294 469958 298350
rect 470014 298294 470082 298350
rect 470138 298294 500678 298350
rect 500734 298294 500802 298350
rect 500858 298294 528970 298350
rect 529026 298294 529094 298350
rect 529150 298294 529218 298350
rect 529274 298294 529342 298350
rect 529398 298294 546970 298350
rect 547026 298294 547094 298350
rect 547150 298294 547218 298350
rect 547274 298294 547342 298350
rect 547398 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 39878 298226
rect 39934 298170 40002 298226
rect 40058 298170 70598 298226
rect 70654 298170 70722 298226
rect 70778 298170 101318 298226
rect 101374 298170 101442 298226
rect 101498 298170 132038 298226
rect 132094 298170 132162 298226
rect 132218 298170 162758 298226
rect 162814 298170 162882 298226
rect 162938 298170 193478 298226
rect 193534 298170 193602 298226
rect 193658 298170 224198 298226
rect 224254 298170 224322 298226
rect 224378 298170 254918 298226
rect 254974 298170 255042 298226
rect 255098 298170 285638 298226
rect 285694 298170 285762 298226
rect 285818 298170 316358 298226
rect 316414 298170 316482 298226
rect 316538 298170 347078 298226
rect 347134 298170 347202 298226
rect 347258 298170 377798 298226
rect 377854 298170 377922 298226
rect 377978 298170 408518 298226
rect 408574 298170 408642 298226
rect 408698 298170 439238 298226
rect 439294 298170 439362 298226
rect 439418 298170 469958 298226
rect 470014 298170 470082 298226
rect 470138 298170 500678 298226
rect 500734 298170 500802 298226
rect 500858 298170 528970 298226
rect 529026 298170 529094 298226
rect 529150 298170 529218 298226
rect 529274 298170 529342 298226
rect 529398 298170 546970 298226
rect 547026 298170 547094 298226
rect 547150 298170 547218 298226
rect 547274 298170 547342 298226
rect 547398 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 39878 298102
rect 39934 298046 40002 298102
rect 40058 298046 70598 298102
rect 70654 298046 70722 298102
rect 70778 298046 101318 298102
rect 101374 298046 101442 298102
rect 101498 298046 132038 298102
rect 132094 298046 132162 298102
rect 132218 298046 162758 298102
rect 162814 298046 162882 298102
rect 162938 298046 193478 298102
rect 193534 298046 193602 298102
rect 193658 298046 224198 298102
rect 224254 298046 224322 298102
rect 224378 298046 254918 298102
rect 254974 298046 255042 298102
rect 255098 298046 285638 298102
rect 285694 298046 285762 298102
rect 285818 298046 316358 298102
rect 316414 298046 316482 298102
rect 316538 298046 347078 298102
rect 347134 298046 347202 298102
rect 347258 298046 377798 298102
rect 377854 298046 377922 298102
rect 377978 298046 408518 298102
rect 408574 298046 408642 298102
rect 408698 298046 439238 298102
rect 439294 298046 439362 298102
rect 439418 298046 469958 298102
rect 470014 298046 470082 298102
rect 470138 298046 500678 298102
rect 500734 298046 500802 298102
rect 500858 298046 528970 298102
rect 529026 298046 529094 298102
rect 529150 298046 529218 298102
rect 529274 298046 529342 298102
rect 529398 298046 546970 298102
rect 547026 298046 547094 298102
rect 547150 298046 547218 298102
rect 547274 298046 547342 298102
rect 547398 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 39878 297978
rect 39934 297922 40002 297978
rect 40058 297922 70598 297978
rect 70654 297922 70722 297978
rect 70778 297922 101318 297978
rect 101374 297922 101442 297978
rect 101498 297922 132038 297978
rect 132094 297922 132162 297978
rect 132218 297922 162758 297978
rect 162814 297922 162882 297978
rect 162938 297922 193478 297978
rect 193534 297922 193602 297978
rect 193658 297922 224198 297978
rect 224254 297922 224322 297978
rect 224378 297922 254918 297978
rect 254974 297922 255042 297978
rect 255098 297922 285638 297978
rect 285694 297922 285762 297978
rect 285818 297922 316358 297978
rect 316414 297922 316482 297978
rect 316538 297922 347078 297978
rect 347134 297922 347202 297978
rect 347258 297922 377798 297978
rect 377854 297922 377922 297978
rect 377978 297922 408518 297978
rect 408574 297922 408642 297978
rect 408698 297922 439238 297978
rect 439294 297922 439362 297978
rect 439418 297922 469958 297978
rect 470014 297922 470082 297978
rect 470138 297922 500678 297978
rect 500734 297922 500802 297978
rect 500858 297922 528970 297978
rect 529026 297922 529094 297978
rect 529150 297922 529218 297978
rect 529274 297922 529342 297978
rect 529398 297922 546970 297978
rect 547026 297922 547094 297978
rect 547150 297922 547218 297978
rect 547274 297922 547342 297978
rect 547398 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 24518 292350
rect 24574 292294 24642 292350
rect 24698 292294 55238 292350
rect 55294 292294 55362 292350
rect 55418 292294 85958 292350
rect 86014 292294 86082 292350
rect 86138 292294 116678 292350
rect 116734 292294 116802 292350
rect 116858 292294 147398 292350
rect 147454 292294 147522 292350
rect 147578 292294 178118 292350
rect 178174 292294 178242 292350
rect 178298 292294 208838 292350
rect 208894 292294 208962 292350
rect 209018 292294 239558 292350
rect 239614 292294 239682 292350
rect 239738 292294 270278 292350
rect 270334 292294 270402 292350
rect 270458 292294 300998 292350
rect 301054 292294 301122 292350
rect 301178 292294 331718 292350
rect 331774 292294 331842 292350
rect 331898 292294 362438 292350
rect 362494 292294 362562 292350
rect 362618 292294 393158 292350
rect 393214 292294 393282 292350
rect 393338 292294 423878 292350
rect 423934 292294 424002 292350
rect 424058 292294 454598 292350
rect 454654 292294 454722 292350
rect 454778 292294 485318 292350
rect 485374 292294 485442 292350
rect 485498 292294 516038 292350
rect 516094 292294 516162 292350
rect 516218 292294 525250 292350
rect 525306 292294 525374 292350
rect 525430 292294 525498 292350
rect 525554 292294 525622 292350
rect 525678 292294 543250 292350
rect 543306 292294 543374 292350
rect 543430 292294 543498 292350
rect 543554 292294 543622 292350
rect 543678 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 24518 292226
rect 24574 292170 24642 292226
rect 24698 292170 55238 292226
rect 55294 292170 55362 292226
rect 55418 292170 85958 292226
rect 86014 292170 86082 292226
rect 86138 292170 116678 292226
rect 116734 292170 116802 292226
rect 116858 292170 147398 292226
rect 147454 292170 147522 292226
rect 147578 292170 178118 292226
rect 178174 292170 178242 292226
rect 178298 292170 208838 292226
rect 208894 292170 208962 292226
rect 209018 292170 239558 292226
rect 239614 292170 239682 292226
rect 239738 292170 270278 292226
rect 270334 292170 270402 292226
rect 270458 292170 300998 292226
rect 301054 292170 301122 292226
rect 301178 292170 331718 292226
rect 331774 292170 331842 292226
rect 331898 292170 362438 292226
rect 362494 292170 362562 292226
rect 362618 292170 393158 292226
rect 393214 292170 393282 292226
rect 393338 292170 423878 292226
rect 423934 292170 424002 292226
rect 424058 292170 454598 292226
rect 454654 292170 454722 292226
rect 454778 292170 485318 292226
rect 485374 292170 485442 292226
rect 485498 292170 516038 292226
rect 516094 292170 516162 292226
rect 516218 292170 525250 292226
rect 525306 292170 525374 292226
rect 525430 292170 525498 292226
rect 525554 292170 525622 292226
rect 525678 292170 543250 292226
rect 543306 292170 543374 292226
rect 543430 292170 543498 292226
rect 543554 292170 543622 292226
rect 543678 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 24518 292102
rect 24574 292046 24642 292102
rect 24698 292046 55238 292102
rect 55294 292046 55362 292102
rect 55418 292046 85958 292102
rect 86014 292046 86082 292102
rect 86138 292046 116678 292102
rect 116734 292046 116802 292102
rect 116858 292046 147398 292102
rect 147454 292046 147522 292102
rect 147578 292046 178118 292102
rect 178174 292046 178242 292102
rect 178298 292046 208838 292102
rect 208894 292046 208962 292102
rect 209018 292046 239558 292102
rect 239614 292046 239682 292102
rect 239738 292046 270278 292102
rect 270334 292046 270402 292102
rect 270458 292046 300998 292102
rect 301054 292046 301122 292102
rect 301178 292046 331718 292102
rect 331774 292046 331842 292102
rect 331898 292046 362438 292102
rect 362494 292046 362562 292102
rect 362618 292046 393158 292102
rect 393214 292046 393282 292102
rect 393338 292046 423878 292102
rect 423934 292046 424002 292102
rect 424058 292046 454598 292102
rect 454654 292046 454722 292102
rect 454778 292046 485318 292102
rect 485374 292046 485442 292102
rect 485498 292046 516038 292102
rect 516094 292046 516162 292102
rect 516218 292046 525250 292102
rect 525306 292046 525374 292102
rect 525430 292046 525498 292102
rect 525554 292046 525622 292102
rect 525678 292046 543250 292102
rect 543306 292046 543374 292102
rect 543430 292046 543498 292102
rect 543554 292046 543622 292102
rect 543678 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 24518 291978
rect 24574 291922 24642 291978
rect 24698 291922 55238 291978
rect 55294 291922 55362 291978
rect 55418 291922 85958 291978
rect 86014 291922 86082 291978
rect 86138 291922 116678 291978
rect 116734 291922 116802 291978
rect 116858 291922 147398 291978
rect 147454 291922 147522 291978
rect 147578 291922 178118 291978
rect 178174 291922 178242 291978
rect 178298 291922 208838 291978
rect 208894 291922 208962 291978
rect 209018 291922 239558 291978
rect 239614 291922 239682 291978
rect 239738 291922 270278 291978
rect 270334 291922 270402 291978
rect 270458 291922 300998 291978
rect 301054 291922 301122 291978
rect 301178 291922 331718 291978
rect 331774 291922 331842 291978
rect 331898 291922 362438 291978
rect 362494 291922 362562 291978
rect 362618 291922 393158 291978
rect 393214 291922 393282 291978
rect 393338 291922 423878 291978
rect 423934 291922 424002 291978
rect 424058 291922 454598 291978
rect 454654 291922 454722 291978
rect 454778 291922 485318 291978
rect 485374 291922 485442 291978
rect 485498 291922 516038 291978
rect 516094 291922 516162 291978
rect 516218 291922 525250 291978
rect 525306 291922 525374 291978
rect 525430 291922 525498 291978
rect 525554 291922 525622 291978
rect 525678 291922 543250 291978
rect 543306 291922 543374 291978
rect 543430 291922 543498 291978
rect 543554 291922 543622 291978
rect 543678 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 39878 280350
rect 39934 280294 40002 280350
rect 40058 280294 70598 280350
rect 70654 280294 70722 280350
rect 70778 280294 101318 280350
rect 101374 280294 101442 280350
rect 101498 280294 132038 280350
rect 132094 280294 132162 280350
rect 132218 280294 162758 280350
rect 162814 280294 162882 280350
rect 162938 280294 193478 280350
rect 193534 280294 193602 280350
rect 193658 280294 224198 280350
rect 224254 280294 224322 280350
rect 224378 280294 254918 280350
rect 254974 280294 255042 280350
rect 255098 280294 285638 280350
rect 285694 280294 285762 280350
rect 285818 280294 316358 280350
rect 316414 280294 316482 280350
rect 316538 280294 347078 280350
rect 347134 280294 347202 280350
rect 347258 280294 377798 280350
rect 377854 280294 377922 280350
rect 377978 280294 408518 280350
rect 408574 280294 408642 280350
rect 408698 280294 439238 280350
rect 439294 280294 439362 280350
rect 439418 280294 469958 280350
rect 470014 280294 470082 280350
rect 470138 280294 500678 280350
rect 500734 280294 500802 280350
rect 500858 280294 528970 280350
rect 529026 280294 529094 280350
rect 529150 280294 529218 280350
rect 529274 280294 529342 280350
rect 529398 280294 546970 280350
rect 547026 280294 547094 280350
rect 547150 280294 547218 280350
rect 547274 280294 547342 280350
rect 547398 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 39878 280226
rect 39934 280170 40002 280226
rect 40058 280170 70598 280226
rect 70654 280170 70722 280226
rect 70778 280170 101318 280226
rect 101374 280170 101442 280226
rect 101498 280170 132038 280226
rect 132094 280170 132162 280226
rect 132218 280170 162758 280226
rect 162814 280170 162882 280226
rect 162938 280170 193478 280226
rect 193534 280170 193602 280226
rect 193658 280170 224198 280226
rect 224254 280170 224322 280226
rect 224378 280170 254918 280226
rect 254974 280170 255042 280226
rect 255098 280170 285638 280226
rect 285694 280170 285762 280226
rect 285818 280170 316358 280226
rect 316414 280170 316482 280226
rect 316538 280170 347078 280226
rect 347134 280170 347202 280226
rect 347258 280170 377798 280226
rect 377854 280170 377922 280226
rect 377978 280170 408518 280226
rect 408574 280170 408642 280226
rect 408698 280170 439238 280226
rect 439294 280170 439362 280226
rect 439418 280170 469958 280226
rect 470014 280170 470082 280226
rect 470138 280170 500678 280226
rect 500734 280170 500802 280226
rect 500858 280170 528970 280226
rect 529026 280170 529094 280226
rect 529150 280170 529218 280226
rect 529274 280170 529342 280226
rect 529398 280170 546970 280226
rect 547026 280170 547094 280226
rect 547150 280170 547218 280226
rect 547274 280170 547342 280226
rect 547398 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 39878 280102
rect 39934 280046 40002 280102
rect 40058 280046 70598 280102
rect 70654 280046 70722 280102
rect 70778 280046 101318 280102
rect 101374 280046 101442 280102
rect 101498 280046 132038 280102
rect 132094 280046 132162 280102
rect 132218 280046 162758 280102
rect 162814 280046 162882 280102
rect 162938 280046 193478 280102
rect 193534 280046 193602 280102
rect 193658 280046 224198 280102
rect 224254 280046 224322 280102
rect 224378 280046 254918 280102
rect 254974 280046 255042 280102
rect 255098 280046 285638 280102
rect 285694 280046 285762 280102
rect 285818 280046 316358 280102
rect 316414 280046 316482 280102
rect 316538 280046 347078 280102
rect 347134 280046 347202 280102
rect 347258 280046 377798 280102
rect 377854 280046 377922 280102
rect 377978 280046 408518 280102
rect 408574 280046 408642 280102
rect 408698 280046 439238 280102
rect 439294 280046 439362 280102
rect 439418 280046 469958 280102
rect 470014 280046 470082 280102
rect 470138 280046 500678 280102
rect 500734 280046 500802 280102
rect 500858 280046 528970 280102
rect 529026 280046 529094 280102
rect 529150 280046 529218 280102
rect 529274 280046 529342 280102
rect 529398 280046 546970 280102
rect 547026 280046 547094 280102
rect 547150 280046 547218 280102
rect 547274 280046 547342 280102
rect 547398 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 39878 279978
rect 39934 279922 40002 279978
rect 40058 279922 70598 279978
rect 70654 279922 70722 279978
rect 70778 279922 101318 279978
rect 101374 279922 101442 279978
rect 101498 279922 132038 279978
rect 132094 279922 132162 279978
rect 132218 279922 162758 279978
rect 162814 279922 162882 279978
rect 162938 279922 193478 279978
rect 193534 279922 193602 279978
rect 193658 279922 224198 279978
rect 224254 279922 224322 279978
rect 224378 279922 254918 279978
rect 254974 279922 255042 279978
rect 255098 279922 285638 279978
rect 285694 279922 285762 279978
rect 285818 279922 316358 279978
rect 316414 279922 316482 279978
rect 316538 279922 347078 279978
rect 347134 279922 347202 279978
rect 347258 279922 377798 279978
rect 377854 279922 377922 279978
rect 377978 279922 408518 279978
rect 408574 279922 408642 279978
rect 408698 279922 439238 279978
rect 439294 279922 439362 279978
rect 439418 279922 469958 279978
rect 470014 279922 470082 279978
rect 470138 279922 500678 279978
rect 500734 279922 500802 279978
rect 500858 279922 528970 279978
rect 529026 279922 529094 279978
rect 529150 279922 529218 279978
rect 529274 279922 529342 279978
rect 529398 279922 546970 279978
rect 547026 279922 547094 279978
rect 547150 279922 547218 279978
rect 547274 279922 547342 279978
rect 547398 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 24518 274350
rect 24574 274294 24642 274350
rect 24698 274294 55238 274350
rect 55294 274294 55362 274350
rect 55418 274294 85958 274350
rect 86014 274294 86082 274350
rect 86138 274294 116678 274350
rect 116734 274294 116802 274350
rect 116858 274294 147398 274350
rect 147454 274294 147522 274350
rect 147578 274294 178118 274350
rect 178174 274294 178242 274350
rect 178298 274294 208838 274350
rect 208894 274294 208962 274350
rect 209018 274294 239558 274350
rect 239614 274294 239682 274350
rect 239738 274294 270278 274350
rect 270334 274294 270402 274350
rect 270458 274294 300998 274350
rect 301054 274294 301122 274350
rect 301178 274294 331718 274350
rect 331774 274294 331842 274350
rect 331898 274294 362438 274350
rect 362494 274294 362562 274350
rect 362618 274294 393158 274350
rect 393214 274294 393282 274350
rect 393338 274294 423878 274350
rect 423934 274294 424002 274350
rect 424058 274294 454598 274350
rect 454654 274294 454722 274350
rect 454778 274294 485318 274350
rect 485374 274294 485442 274350
rect 485498 274294 516038 274350
rect 516094 274294 516162 274350
rect 516218 274294 525250 274350
rect 525306 274294 525374 274350
rect 525430 274294 525498 274350
rect 525554 274294 525622 274350
rect 525678 274294 543250 274350
rect 543306 274294 543374 274350
rect 543430 274294 543498 274350
rect 543554 274294 543622 274350
rect 543678 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 24518 274226
rect 24574 274170 24642 274226
rect 24698 274170 55238 274226
rect 55294 274170 55362 274226
rect 55418 274170 85958 274226
rect 86014 274170 86082 274226
rect 86138 274170 116678 274226
rect 116734 274170 116802 274226
rect 116858 274170 147398 274226
rect 147454 274170 147522 274226
rect 147578 274170 178118 274226
rect 178174 274170 178242 274226
rect 178298 274170 208838 274226
rect 208894 274170 208962 274226
rect 209018 274170 239558 274226
rect 239614 274170 239682 274226
rect 239738 274170 270278 274226
rect 270334 274170 270402 274226
rect 270458 274170 300998 274226
rect 301054 274170 301122 274226
rect 301178 274170 331718 274226
rect 331774 274170 331842 274226
rect 331898 274170 362438 274226
rect 362494 274170 362562 274226
rect 362618 274170 393158 274226
rect 393214 274170 393282 274226
rect 393338 274170 423878 274226
rect 423934 274170 424002 274226
rect 424058 274170 454598 274226
rect 454654 274170 454722 274226
rect 454778 274170 485318 274226
rect 485374 274170 485442 274226
rect 485498 274170 516038 274226
rect 516094 274170 516162 274226
rect 516218 274170 525250 274226
rect 525306 274170 525374 274226
rect 525430 274170 525498 274226
rect 525554 274170 525622 274226
rect 525678 274170 543250 274226
rect 543306 274170 543374 274226
rect 543430 274170 543498 274226
rect 543554 274170 543622 274226
rect 543678 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 24518 274102
rect 24574 274046 24642 274102
rect 24698 274046 55238 274102
rect 55294 274046 55362 274102
rect 55418 274046 85958 274102
rect 86014 274046 86082 274102
rect 86138 274046 116678 274102
rect 116734 274046 116802 274102
rect 116858 274046 147398 274102
rect 147454 274046 147522 274102
rect 147578 274046 178118 274102
rect 178174 274046 178242 274102
rect 178298 274046 208838 274102
rect 208894 274046 208962 274102
rect 209018 274046 239558 274102
rect 239614 274046 239682 274102
rect 239738 274046 270278 274102
rect 270334 274046 270402 274102
rect 270458 274046 300998 274102
rect 301054 274046 301122 274102
rect 301178 274046 331718 274102
rect 331774 274046 331842 274102
rect 331898 274046 362438 274102
rect 362494 274046 362562 274102
rect 362618 274046 393158 274102
rect 393214 274046 393282 274102
rect 393338 274046 423878 274102
rect 423934 274046 424002 274102
rect 424058 274046 454598 274102
rect 454654 274046 454722 274102
rect 454778 274046 485318 274102
rect 485374 274046 485442 274102
rect 485498 274046 516038 274102
rect 516094 274046 516162 274102
rect 516218 274046 525250 274102
rect 525306 274046 525374 274102
rect 525430 274046 525498 274102
rect 525554 274046 525622 274102
rect 525678 274046 543250 274102
rect 543306 274046 543374 274102
rect 543430 274046 543498 274102
rect 543554 274046 543622 274102
rect 543678 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 24518 273978
rect 24574 273922 24642 273978
rect 24698 273922 55238 273978
rect 55294 273922 55362 273978
rect 55418 273922 85958 273978
rect 86014 273922 86082 273978
rect 86138 273922 116678 273978
rect 116734 273922 116802 273978
rect 116858 273922 147398 273978
rect 147454 273922 147522 273978
rect 147578 273922 178118 273978
rect 178174 273922 178242 273978
rect 178298 273922 208838 273978
rect 208894 273922 208962 273978
rect 209018 273922 239558 273978
rect 239614 273922 239682 273978
rect 239738 273922 270278 273978
rect 270334 273922 270402 273978
rect 270458 273922 300998 273978
rect 301054 273922 301122 273978
rect 301178 273922 331718 273978
rect 331774 273922 331842 273978
rect 331898 273922 362438 273978
rect 362494 273922 362562 273978
rect 362618 273922 393158 273978
rect 393214 273922 393282 273978
rect 393338 273922 423878 273978
rect 423934 273922 424002 273978
rect 424058 273922 454598 273978
rect 454654 273922 454722 273978
rect 454778 273922 485318 273978
rect 485374 273922 485442 273978
rect 485498 273922 516038 273978
rect 516094 273922 516162 273978
rect 516218 273922 525250 273978
rect 525306 273922 525374 273978
rect 525430 273922 525498 273978
rect 525554 273922 525622 273978
rect 525678 273922 543250 273978
rect 543306 273922 543374 273978
rect 543430 273922 543498 273978
rect 543554 273922 543622 273978
rect 543678 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 39878 262350
rect 39934 262294 40002 262350
rect 40058 262294 70598 262350
rect 70654 262294 70722 262350
rect 70778 262294 101318 262350
rect 101374 262294 101442 262350
rect 101498 262294 132038 262350
rect 132094 262294 132162 262350
rect 132218 262294 162758 262350
rect 162814 262294 162882 262350
rect 162938 262294 193478 262350
rect 193534 262294 193602 262350
rect 193658 262294 224198 262350
rect 224254 262294 224322 262350
rect 224378 262294 254918 262350
rect 254974 262294 255042 262350
rect 255098 262294 285638 262350
rect 285694 262294 285762 262350
rect 285818 262294 316358 262350
rect 316414 262294 316482 262350
rect 316538 262294 347078 262350
rect 347134 262294 347202 262350
rect 347258 262294 377798 262350
rect 377854 262294 377922 262350
rect 377978 262294 408518 262350
rect 408574 262294 408642 262350
rect 408698 262294 439238 262350
rect 439294 262294 439362 262350
rect 439418 262294 469958 262350
rect 470014 262294 470082 262350
rect 470138 262294 500678 262350
rect 500734 262294 500802 262350
rect 500858 262294 528970 262350
rect 529026 262294 529094 262350
rect 529150 262294 529218 262350
rect 529274 262294 529342 262350
rect 529398 262294 546970 262350
rect 547026 262294 547094 262350
rect 547150 262294 547218 262350
rect 547274 262294 547342 262350
rect 547398 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 39878 262226
rect 39934 262170 40002 262226
rect 40058 262170 70598 262226
rect 70654 262170 70722 262226
rect 70778 262170 101318 262226
rect 101374 262170 101442 262226
rect 101498 262170 132038 262226
rect 132094 262170 132162 262226
rect 132218 262170 162758 262226
rect 162814 262170 162882 262226
rect 162938 262170 193478 262226
rect 193534 262170 193602 262226
rect 193658 262170 224198 262226
rect 224254 262170 224322 262226
rect 224378 262170 254918 262226
rect 254974 262170 255042 262226
rect 255098 262170 285638 262226
rect 285694 262170 285762 262226
rect 285818 262170 316358 262226
rect 316414 262170 316482 262226
rect 316538 262170 347078 262226
rect 347134 262170 347202 262226
rect 347258 262170 377798 262226
rect 377854 262170 377922 262226
rect 377978 262170 408518 262226
rect 408574 262170 408642 262226
rect 408698 262170 439238 262226
rect 439294 262170 439362 262226
rect 439418 262170 469958 262226
rect 470014 262170 470082 262226
rect 470138 262170 500678 262226
rect 500734 262170 500802 262226
rect 500858 262170 528970 262226
rect 529026 262170 529094 262226
rect 529150 262170 529218 262226
rect 529274 262170 529342 262226
rect 529398 262170 546970 262226
rect 547026 262170 547094 262226
rect 547150 262170 547218 262226
rect 547274 262170 547342 262226
rect 547398 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 39878 262102
rect 39934 262046 40002 262102
rect 40058 262046 70598 262102
rect 70654 262046 70722 262102
rect 70778 262046 101318 262102
rect 101374 262046 101442 262102
rect 101498 262046 132038 262102
rect 132094 262046 132162 262102
rect 132218 262046 162758 262102
rect 162814 262046 162882 262102
rect 162938 262046 193478 262102
rect 193534 262046 193602 262102
rect 193658 262046 224198 262102
rect 224254 262046 224322 262102
rect 224378 262046 254918 262102
rect 254974 262046 255042 262102
rect 255098 262046 285638 262102
rect 285694 262046 285762 262102
rect 285818 262046 316358 262102
rect 316414 262046 316482 262102
rect 316538 262046 347078 262102
rect 347134 262046 347202 262102
rect 347258 262046 377798 262102
rect 377854 262046 377922 262102
rect 377978 262046 408518 262102
rect 408574 262046 408642 262102
rect 408698 262046 439238 262102
rect 439294 262046 439362 262102
rect 439418 262046 469958 262102
rect 470014 262046 470082 262102
rect 470138 262046 500678 262102
rect 500734 262046 500802 262102
rect 500858 262046 528970 262102
rect 529026 262046 529094 262102
rect 529150 262046 529218 262102
rect 529274 262046 529342 262102
rect 529398 262046 546970 262102
rect 547026 262046 547094 262102
rect 547150 262046 547218 262102
rect 547274 262046 547342 262102
rect 547398 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 39878 261978
rect 39934 261922 40002 261978
rect 40058 261922 70598 261978
rect 70654 261922 70722 261978
rect 70778 261922 101318 261978
rect 101374 261922 101442 261978
rect 101498 261922 132038 261978
rect 132094 261922 132162 261978
rect 132218 261922 162758 261978
rect 162814 261922 162882 261978
rect 162938 261922 193478 261978
rect 193534 261922 193602 261978
rect 193658 261922 224198 261978
rect 224254 261922 224322 261978
rect 224378 261922 254918 261978
rect 254974 261922 255042 261978
rect 255098 261922 285638 261978
rect 285694 261922 285762 261978
rect 285818 261922 316358 261978
rect 316414 261922 316482 261978
rect 316538 261922 347078 261978
rect 347134 261922 347202 261978
rect 347258 261922 377798 261978
rect 377854 261922 377922 261978
rect 377978 261922 408518 261978
rect 408574 261922 408642 261978
rect 408698 261922 439238 261978
rect 439294 261922 439362 261978
rect 439418 261922 469958 261978
rect 470014 261922 470082 261978
rect 470138 261922 500678 261978
rect 500734 261922 500802 261978
rect 500858 261922 528970 261978
rect 529026 261922 529094 261978
rect 529150 261922 529218 261978
rect 529274 261922 529342 261978
rect 529398 261922 546970 261978
rect 547026 261922 547094 261978
rect 547150 261922 547218 261978
rect 547274 261922 547342 261978
rect 547398 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 24518 256350
rect 24574 256294 24642 256350
rect 24698 256294 55238 256350
rect 55294 256294 55362 256350
rect 55418 256294 85958 256350
rect 86014 256294 86082 256350
rect 86138 256294 116678 256350
rect 116734 256294 116802 256350
rect 116858 256294 147398 256350
rect 147454 256294 147522 256350
rect 147578 256294 178118 256350
rect 178174 256294 178242 256350
rect 178298 256294 208838 256350
rect 208894 256294 208962 256350
rect 209018 256294 239558 256350
rect 239614 256294 239682 256350
rect 239738 256294 270278 256350
rect 270334 256294 270402 256350
rect 270458 256294 300998 256350
rect 301054 256294 301122 256350
rect 301178 256294 331718 256350
rect 331774 256294 331842 256350
rect 331898 256294 362438 256350
rect 362494 256294 362562 256350
rect 362618 256294 393158 256350
rect 393214 256294 393282 256350
rect 393338 256294 423878 256350
rect 423934 256294 424002 256350
rect 424058 256294 454598 256350
rect 454654 256294 454722 256350
rect 454778 256294 485318 256350
rect 485374 256294 485442 256350
rect 485498 256294 516038 256350
rect 516094 256294 516162 256350
rect 516218 256294 525250 256350
rect 525306 256294 525374 256350
rect 525430 256294 525498 256350
rect 525554 256294 525622 256350
rect 525678 256294 543250 256350
rect 543306 256294 543374 256350
rect 543430 256294 543498 256350
rect 543554 256294 543622 256350
rect 543678 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 24518 256226
rect 24574 256170 24642 256226
rect 24698 256170 55238 256226
rect 55294 256170 55362 256226
rect 55418 256170 85958 256226
rect 86014 256170 86082 256226
rect 86138 256170 116678 256226
rect 116734 256170 116802 256226
rect 116858 256170 147398 256226
rect 147454 256170 147522 256226
rect 147578 256170 178118 256226
rect 178174 256170 178242 256226
rect 178298 256170 208838 256226
rect 208894 256170 208962 256226
rect 209018 256170 239558 256226
rect 239614 256170 239682 256226
rect 239738 256170 270278 256226
rect 270334 256170 270402 256226
rect 270458 256170 300998 256226
rect 301054 256170 301122 256226
rect 301178 256170 331718 256226
rect 331774 256170 331842 256226
rect 331898 256170 362438 256226
rect 362494 256170 362562 256226
rect 362618 256170 393158 256226
rect 393214 256170 393282 256226
rect 393338 256170 423878 256226
rect 423934 256170 424002 256226
rect 424058 256170 454598 256226
rect 454654 256170 454722 256226
rect 454778 256170 485318 256226
rect 485374 256170 485442 256226
rect 485498 256170 516038 256226
rect 516094 256170 516162 256226
rect 516218 256170 525250 256226
rect 525306 256170 525374 256226
rect 525430 256170 525498 256226
rect 525554 256170 525622 256226
rect 525678 256170 543250 256226
rect 543306 256170 543374 256226
rect 543430 256170 543498 256226
rect 543554 256170 543622 256226
rect 543678 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 24518 256102
rect 24574 256046 24642 256102
rect 24698 256046 55238 256102
rect 55294 256046 55362 256102
rect 55418 256046 85958 256102
rect 86014 256046 86082 256102
rect 86138 256046 116678 256102
rect 116734 256046 116802 256102
rect 116858 256046 147398 256102
rect 147454 256046 147522 256102
rect 147578 256046 178118 256102
rect 178174 256046 178242 256102
rect 178298 256046 208838 256102
rect 208894 256046 208962 256102
rect 209018 256046 239558 256102
rect 239614 256046 239682 256102
rect 239738 256046 270278 256102
rect 270334 256046 270402 256102
rect 270458 256046 300998 256102
rect 301054 256046 301122 256102
rect 301178 256046 331718 256102
rect 331774 256046 331842 256102
rect 331898 256046 362438 256102
rect 362494 256046 362562 256102
rect 362618 256046 393158 256102
rect 393214 256046 393282 256102
rect 393338 256046 423878 256102
rect 423934 256046 424002 256102
rect 424058 256046 454598 256102
rect 454654 256046 454722 256102
rect 454778 256046 485318 256102
rect 485374 256046 485442 256102
rect 485498 256046 516038 256102
rect 516094 256046 516162 256102
rect 516218 256046 525250 256102
rect 525306 256046 525374 256102
rect 525430 256046 525498 256102
rect 525554 256046 525622 256102
rect 525678 256046 543250 256102
rect 543306 256046 543374 256102
rect 543430 256046 543498 256102
rect 543554 256046 543622 256102
rect 543678 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 24518 255978
rect 24574 255922 24642 255978
rect 24698 255922 55238 255978
rect 55294 255922 55362 255978
rect 55418 255922 85958 255978
rect 86014 255922 86082 255978
rect 86138 255922 116678 255978
rect 116734 255922 116802 255978
rect 116858 255922 147398 255978
rect 147454 255922 147522 255978
rect 147578 255922 178118 255978
rect 178174 255922 178242 255978
rect 178298 255922 208838 255978
rect 208894 255922 208962 255978
rect 209018 255922 239558 255978
rect 239614 255922 239682 255978
rect 239738 255922 270278 255978
rect 270334 255922 270402 255978
rect 270458 255922 300998 255978
rect 301054 255922 301122 255978
rect 301178 255922 331718 255978
rect 331774 255922 331842 255978
rect 331898 255922 362438 255978
rect 362494 255922 362562 255978
rect 362618 255922 393158 255978
rect 393214 255922 393282 255978
rect 393338 255922 423878 255978
rect 423934 255922 424002 255978
rect 424058 255922 454598 255978
rect 454654 255922 454722 255978
rect 454778 255922 485318 255978
rect 485374 255922 485442 255978
rect 485498 255922 516038 255978
rect 516094 255922 516162 255978
rect 516218 255922 525250 255978
rect 525306 255922 525374 255978
rect 525430 255922 525498 255978
rect 525554 255922 525622 255978
rect 525678 255922 543250 255978
rect 543306 255922 543374 255978
rect 543430 255922 543498 255978
rect 543554 255922 543622 255978
rect 543678 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 39878 244350
rect 39934 244294 40002 244350
rect 40058 244294 70598 244350
rect 70654 244294 70722 244350
rect 70778 244294 101318 244350
rect 101374 244294 101442 244350
rect 101498 244294 132038 244350
rect 132094 244294 132162 244350
rect 132218 244294 162758 244350
rect 162814 244294 162882 244350
rect 162938 244294 193478 244350
rect 193534 244294 193602 244350
rect 193658 244294 224198 244350
rect 224254 244294 224322 244350
rect 224378 244294 254918 244350
rect 254974 244294 255042 244350
rect 255098 244294 285638 244350
rect 285694 244294 285762 244350
rect 285818 244294 316358 244350
rect 316414 244294 316482 244350
rect 316538 244294 347078 244350
rect 347134 244294 347202 244350
rect 347258 244294 377798 244350
rect 377854 244294 377922 244350
rect 377978 244294 408518 244350
rect 408574 244294 408642 244350
rect 408698 244294 439238 244350
rect 439294 244294 439362 244350
rect 439418 244294 469958 244350
rect 470014 244294 470082 244350
rect 470138 244294 500678 244350
rect 500734 244294 500802 244350
rect 500858 244294 528970 244350
rect 529026 244294 529094 244350
rect 529150 244294 529218 244350
rect 529274 244294 529342 244350
rect 529398 244294 546970 244350
rect 547026 244294 547094 244350
rect 547150 244294 547218 244350
rect 547274 244294 547342 244350
rect 547398 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 39878 244226
rect 39934 244170 40002 244226
rect 40058 244170 70598 244226
rect 70654 244170 70722 244226
rect 70778 244170 101318 244226
rect 101374 244170 101442 244226
rect 101498 244170 132038 244226
rect 132094 244170 132162 244226
rect 132218 244170 162758 244226
rect 162814 244170 162882 244226
rect 162938 244170 193478 244226
rect 193534 244170 193602 244226
rect 193658 244170 224198 244226
rect 224254 244170 224322 244226
rect 224378 244170 254918 244226
rect 254974 244170 255042 244226
rect 255098 244170 285638 244226
rect 285694 244170 285762 244226
rect 285818 244170 316358 244226
rect 316414 244170 316482 244226
rect 316538 244170 347078 244226
rect 347134 244170 347202 244226
rect 347258 244170 377798 244226
rect 377854 244170 377922 244226
rect 377978 244170 408518 244226
rect 408574 244170 408642 244226
rect 408698 244170 439238 244226
rect 439294 244170 439362 244226
rect 439418 244170 469958 244226
rect 470014 244170 470082 244226
rect 470138 244170 500678 244226
rect 500734 244170 500802 244226
rect 500858 244170 528970 244226
rect 529026 244170 529094 244226
rect 529150 244170 529218 244226
rect 529274 244170 529342 244226
rect 529398 244170 546970 244226
rect 547026 244170 547094 244226
rect 547150 244170 547218 244226
rect 547274 244170 547342 244226
rect 547398 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 39878 244102
rect 39934 244046 40002 244102
rect 40058 244046 70598 244102
rect 70654 244046 70722 244102
rect 70778 244046 101318 244102
rect 101374 244046 101442 244102
rect 101498 244046 132038 244102
rect 132094 244046 132162 244102
rect 132218 244046 162758 244102
rect 162814 244046 162882 244102
rect 162938 244046 193478 244102
rect 193534 244046 193602 244102
rect 193658 244046 224198 244102
rect 224254 244046 224322 244102
rect 224378 244046 254918 244102
rect 254974 244046 255042 244102
rect 255098 244046 285638 244102
rect 285694 244046 285762 244102
rect 285818 244046 316358 244102
rect 316414 244046 316482 244102
rect 316538 244046 347078 244102
rect 347134 244046 347202 244102
rect 347258 244046 377798 244102
rect 377854 244046 377922 244102
rect 377978 244046 408518 244102
rect 408574 244046 408642 244102
rect 408698 244046 439238 244102
rect 439294 244046 439362 244102
rect 439418 244046 469958 244102
rect 470014 244046 470082 244102
rect 470138 244046 500678 244102
rect 500734 244046 500802 244102
rect 500858 244046 528970 244102
rect 529026 244046 529094 244102
rect 529150 244046 529218 244102
rect 529274 244046 529342 244102
rect 529398 244046 546970 244102
rect 547026 244046 547094 244102
rect 547150 244046 547218 244102
rect 547274 244046 547342 244102
rect 547398 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 39878 243978
rect 39934 243922 40002 243978
rect 40058 243922 70598 243978
rect 70654 243922 70722 243978
rect 70778 243922 101318 243978
rect 101374 243922 101442 243978
rect 101498 243922 132038 243978
rect 132094 243922 132162 243978
rect 132218 243922 162758 243978
rect 162814 243922 162882 243978
rect 162938 243922 193478 243978
rect 193534 243922 193602 243978
rect 193658 243922 224198 243978
rect 224254 243922 224322 243978
rect 224378 243922 254918 243978
rect 254974 243922 255042 243978
rect 255098 243922 285638 243978
rect 285694 243922 285762 243978
rect 285818 243922 316358 243978
rect 316414 243922 316482 243978
rect 316538 243922 347078 243978
rect 347134 243922 347202 243978
rect 347258 243922 377798 243978
rect 377854 243922 377922 243978
rect 377978 243922 408518 243978
rect 408574 243922 408642 243978
rect 408698 243922 439238 243978
rect 439294 243922 439362 243978
rect 439418 243922 469958 243978
rect 470014 243922 470082 243978
rect 470138 243922 500678 243978
rect 500734 243922 500802 243978
rect 500858 243922 528970 243978
rect 529026 243922 529094 243978
rect 529150 243922 529218 243978
rect 529274 243922 529342 243978
rect 529398 243922 546970 243978
rect 547026 243922 547094 243978
rect 547150 243922 547218 243978
rect 547274 243922 547342 243978
rect 547398 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 24518 238350
rect 24574 238294 24642 238350
rect 24698 238294 55238 238350
rect 55294 238294 55362 238350
rect 55418 238294 85958 238350
rect 86014 238294 86082 238350
rect 86138 238294 116678 238350
rect 116734 238294 116802 238350
rect 116858 238294 147398 238350
rect 147454 238294 147522 238350
rect 147578 238294 178118 238350
rect 178174 238294 178242 238350
rect 178298 238294 208838 238350
rect 208894 238294 208962 238350
rect 209018 238294 239558 238350
rect 239614 238294 239682 238350
rect 239738 238294 270278 238350
rect 270334 238294 270402 238350
rect 270458 238294 300998 238350
rect 301054 238294 301122 238350
rect 301178 238294 331718 238350
rect 331774 238294 331842 238350
rect 331898 238294 362438 238350
rect 362494 238294 362562 238350
rect 362618 238294 393158 238350
rect 393214 238294 393282 238350
rect 393338 238294 423878 238350
rect 423934 238294 424002 238350
rect 424058 238294 454598 238350
rect 454654 238294 454722 238350
rect 454778 238294 485318 238350
rect 485374 238294 485442 238350
rect 485498 238294 516038 238350
rect 516094 238294 516162 238350
rect 516218 238294 525250 238350
rect 525306 238294 525374 238350
rect 525430 238294 525498 238350
rect 525554 238294 525622 238350
rect 525678 238294 543250 238350
rect 543306 238294 543374 238350
rect 543430 238294 543498 238350
rect 543554 238294 543622 238350
rect 543678 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 24518 238226
rect 24574 238170 24642 238226
rect 24698 238170 55238 238226
rect 55294 238170 55362 238226
rect 55418 238170 85958 238226
rect 86014 238170 86082 238226
rect 86138 238170 116678 238226
rect 116734 238170 116802 238226
rect 116858 238170 147398 238226
rect 147454 238170 147522 238226
rect 147578 238170 178118 238226
rect 178174 238170 178242 238226
rect 178298 238170 208838 238226
rect 208894 238170 208962 238226
rect 209018 238170 239558 238226
rect 239614 238170 239682 238226
rect 239738 238170 270278 238226
rect 270334 238170 270402 238226
rect 270458 238170 300998 238226
rect 301054 238170 301122 238226
rect 301178 238170 331718 238226
rect 331774 238170 331842 238226
rect 331898 238170 362438 238226
rect 362494 238170 362562 238226
rect 362618 238170 393158 238226
rect 393214 238170 393282 238226
rect 393338 238170 423878 238226
rect 423934 238170 424002 238226
rect 424058 238170 454598 238226
rect 454654 238170 454722 238226
rect 454778 238170 485318 238226
rect 485374 238170 485442 238226
rect 485498 238170 516038 238226
rect 516094 238170 516162 238226
rect 516218 238170 525250 238226
rect 525306 238170 525374 238226
rect 525430 238170 525498 238226
rect 525554 238170 525622 238226
rect 525678 238170 543250 238226
rect 543306 238170 543374 238226
rect 543430 238170 543498 238226
rect 543554 238170 543622 238226
rect 543678 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 24518 238102
rect 24574 238046 24642 238102
rect 24698 238046 55238 238102
rect 55294 238046 55362 238102
rect 55418 238046 85958 238102
rect 86014 238046 86082 238102
rect 86138 238046 116678 238102
rect 116734 238046 116802 238102
rect 116858 238046 147398 238102
rect 147454 238046 147522 238102
rect 147578 238046 178118 238102
rect 178174 238046 178242 238102
rect 178298 238046 208838 238102
rect 208894 238046 208962 238102
rect 209018 238046 239558 238102
rect 239614 238046 239682 238102
rect 239738 238046 270278 238102
rect 270334 238046 270402 238102
rect 270458 238046 300998 238102
rect 301054 238046 301122 238102
rect 301178 238046 331718 238102
rect 331774 238046 331842 238102
rect 331898 238046 362438 238102
rect 362494 238046 362562 238102
rect 362618 238046 393158 238102
rect 393214 238046 393282 238102
rect 393338 238046 423878 238102
rect 423934 238046 424002 238102
rect 424058 238046 454598 238102
rect 454654 238046 454722 238102
rect 454778 238046 485318 238102
rect 485374 238046 485442 238102
rect 485498 238046 516038 238102
rect 516094 238046 516162 238102
rect 516218 238046 525250 238102
rect 525306 238046 525374 238102
rect 525430 238046 525498 238102
rect 525554 238046 525622 238102
rect 525678 238046 543250 238102
rect 543306 238046 543374 238102
rect 543430 238046 543498 238102
rect 543554 238046 543622 238102
rect 543678 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 24518 237978
rect 24574 237922 24642 237978
rect 24698 237922 55238 237978
rect 55294 237922 55362 237978
rect 55418 237922 85958 237978
rect 86014 237922 86082 237978
rect 86138 237922 116678 237978
rect 116734 237922 116802 237978
rect 116858 237922 147398 237978
rect 147454 237922 147522 237978
rect 147578 237922 178118 237978
rect 178174 237922 178242 237978
rect 178298 237922 208838 237978
rect 208894 237922 208962 237978
rect 209018 237922 239558 237978
rect 239614 237922 239682 237978
rect 239738 237922 270278 237978
rect 270334 237922 270402 237978
rect 270458 237922 300998 237978
rect 301054 237922 301122 237978
rect 301178 237922 331718 237978
rect 331774 237922 331842 237978
rect 331898 237922 362438 237978
rect 362494 237922 362562 237978
rect 362618 237922 393158 237978
rect 393214 237922 393282 237978
rect 393338 237922 423878 237978
rect 423934 237922 424002 237978
rect 424058 237922 454598 237978
rect 454654 237922 454722 237978
rect 454778 237922 485318 237978
rect 485374 237922 485442 237978
rect 485498 237922 516038 237978
rect 516094 237922 516162 237978
rect 516218 237922 525250 237978
rect 525306 237922 525374 237978
rect 525430 237922 525498 237978
rect 525554 237922 525622 237978
rect 525678 237922 543250 237978
rect 543306 237922 543374 237978
rect 543430 237922 543498 237978
rect 543554 237922 543622 237978
rect 543678 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 39878 226350
rect 39934 226294 40002 226350
rect 40058 226294 70598 226350
rect 70654 226294 70722 226350
rect 70778 226294 101318 226350
rect 101374 226294 101442 226350
rect 101498 226294 132038 226350
rect 132094 226294 132162 226350
rect 132218 226294 162758 226350
rect 162814 226294 162882 226350
rect 162938 226294 193478 226350
rect 193534 226294 193602 226350
rect 193658 226294 224198 226350
rect 224254 226294 224322 226350
rect 224378 226294 254918 226350
rect 254974 226294 255042 226350
rect 255098 226294 285638 226350
rect 285694 226294 285762 226350
rect 285818 226294 316358 226350
rect 316414 226294 316482 226350
rect 316538 226294 347078 226350
rect 347134 226294 347202 226350
rect 347258 226294 377798 226350
rect 377854 226294 377922 226350
rect 377978 226294 408518 226350
rect 408574 226294 408642 226350
rect 408698 226294 439238 226350
rect 439294 226294 439362 226350
rect 439418 226294 469958 226350
rect 470014 226294 470082 226350
rect 470138 226294 500678 226350
rect 500734 226294 500802 226350
rect 500858 226294 528970 226350
rect 529026 226294 529094 226350
rect 529150 226294 529218 226350
rect 529274 226294 529342 226350
rect 529398 226294 546970 226350
rect 547026 226294 547094 226350
rect 547150 226294 547218 226350
rect 547274 226294 547342 226350
rect 547398 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 39878 226226
rect 39934 226170 40002 226226
rect 40058 226170 70598 226226
rect 70654 226170 70722 226226
rect 70778 226170 101318 226226
rect 101374 226170 101442 226226
rect 101498 226170 132038 226226
rect 132094 226170 132162 226226
rect 132218 226170 162758 226226
rect 162814 226170 162882 226226
rect 162938 226170 193478 226226
rect 193534 226170 193602 226226
rect 193658 226170 224198 226226
rect 224254 226170 224322 226226
rect 224378 226170 254918 226226
rect 254974 226170 255042 226226
rect 255098 226170 285638 226226
rect 285694 226170 285762 226226
rect 285818 226170 316358 226226
rect 316414 226170 316482 226226
rect 316538 226170 347078 226226
rect 347134 226170 347202 226226
rect 347258 226170 377798 226226
rect 377854 226170 377922 226226
rect 377978 226170 408518 226226
rect 408574 226170 408642 226226
rect 408698 226170 439238 226226
rect 439294 226170 439362 226226
rect 439418 226170 469958 226226
rect 470014 226170 470082 226226
rect 470138 226170 500678 226226
rect 500734 226170 500802 226226
rect 500858 226170 528970 226226
rect 529026 226170 529094 226226
rect 529150 226170 529218 226226
rect 529274 226170 529342 226226
rect 529398 226170 546970 226226
rect 547026 226170 547094 226226
rect 547150 226170 547218 226226
rect 547274 226170 547342 226226
rect 547398 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 39878 226102
rect 39934 226046 40002 226102
rect 40058 226046 70598 226102
rect 70654 226046 70722 226102
rect 70778 226046 101318 226102
rect 101374 226046 101442 226102
rect 101498 226046 132038 226102
rect 132094 226046 132162 226102
rect 132218 226046 162758 226102
rect 162814 226046 162882 226102
rect 162938 226046 193478 226102
rect 193534 226046 193602 226102
rect 193658 226046 224198 226102
rect 224254 226046 224322 226102
rect 224378 226046 254918 226102
rect 254974 226046 255042 226102
rect 255098 226046 285638 226102
rect 285694 226046 285762 226102
rect 285818 226046 316358 226102
rect 316414 226046 316482 226102
rect 316538 226046 347078 226102
rect 347134 226046 347202 226102
rect 347258 226046 377798 226102
rect 377854 226046 377922 226102
rect 377978 226046 408518 226102
rect 408574 226046 408642 226102
rect 408698 226046 439238 226102
rect 439294 226046 439362 226102
rect 439418 226046 469958 226102
rect 470014 226046 470082 226102
rect 470138 226046 500678 226102
rect 500734 226046 500802 226102
rect 500858 226046 528970 226102
rect 529026 226046 529094 226102
rect 529150 226046 529218 226102
rect 529274 226046 529342 226102
rect 529398 226046 546970 226102
rect 547026 226046 547094 226102
rect 547150 226046 547218 226102
rect 547274 226046 547342 226102
rect 547398 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 39878 225978
rect 39934 225922 40002 225978
rect 40058 225922 70598 225978
rect 70654 225922 70722 225978
rect 70778 225922 101318 225978
rect 101374 225922 101442 225978
rect 101498 225922 132038 225978
rect 132094 225922 132162 225978
rect 132218 225922 162758 225978
rect 162814 225922 162882 225978
rect 162938 225922 193478 225978
rect 193534 225922 193602 225978
rect 193658 225922 224198 225978
rect 224254 225922 224322 225978
rect 224378 225922 254918 225978
rect 254974 225922 255042 225978
rect 255098 225922 285638 225978
rect 285694 225922 285762 225978
rect 285818 225922 316358 225978
rect 316414 225922 316482 225978
rect 316538 225922 347078 225978
rect 347134 225922 347202 225978
rect 347258 225922 377798 225978
rect 377854 225922 377922 225978
rect 377978 225922 408518 225978
rect 408574 225922 408642 225978
rect 408698 225922 439238 225978
rect 439294 225922 439362 225978
rect 439418 225922 469958 225978
rect 470014 225922 470082 225978
rect 470138 225922 500678 225978
rect 500734 225922 500802 225978
rect 500858 225922 528970 225978
rect 529026 225922 529094 225978
rect 529150 225922 529218 225978
rect 529274 225922 529342 225978
rect 529398 225922 546970 225978
rect 547026 225922 547094 225978
rect 547150 225922 547218 225978
rect 547274 225922 547342 225978
rect 547398 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 24518 220350
rect 24574 220294 24642 220350
rect 24698 220294 55238 220350
rect 55294 220294 55362 220350
rect 55418 220294 85958 220350
rect 86014 220294 86082 220350
rect 86138 220294 116678 220350
rect 116734 220294 116802 220350
rect 116858 220294 147398 220350
rect 147454 220294 147522 220350
rect 147578 220294 178118 220350
rect 178174 220294 178242 220350
rect 178298 220294 208838 220350
rect 208894 220294 208962 220350
rect 209018 220294 239558 220350
rect 239614 220294 239682 220350
rect 239738 220294 270278 220350
rect 270334 220294 270402 220350
rect 270458 220294 300998 220350
rect 301054 220294 301122 220350
rect 301178 220294 331718 220350
rect 331774 220294 331842 220350
rect 331898 220294 362438 220350
rect 362494 220294 362562 220350
rect 362618 220294 393158 220350
rect 393214 220294 393282 220350
rect 393338 220294 423878 220350
rect 423934 220294 424002 220350
rect 424058 220294 454598 220350
rect 454654 220294 454722 220350
rect 454778 220294 485318 220350
rect 485374 220294 485442 220350
rect 485498 220294 516038 220350
rect 516094 220294 516162 220350
rect 516218 220294 525250 220350
rect 525306 220294 525374 220350
rect 525430 220294 525498 220350
rect 525554 220294 525622 220350
rect 525678 220294 543250 220350
rect 543306 220294 543374 220350
rect 543430 220294 543498 220350
rect 543554 220294 543622 220350
rect 543678 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 24518 220226
rect 24574 220170 24642 220226
rect 24698 220170 55238 220226
rect 55294 220170 55362 220226
rect 55418 220170 85958 220226
rect 86014 220170 86082 220226
rect 86138 220170 116678 220226
rect 116734 220170 116802 220226
rect 116858 220170 147398 220226
rect 147454 220170 147522 220226
rect 147578 220170 178118 220226
rect 178174 220170 178242 220226
rect 178298 220170 208838 220226
rect 208894 220170 208962 220226
rect 209018 220170 239558 220226
rect 239614 220170 239682 220226
rect 239738 220170 270278 220226
rect 270334 220170 270402 220226
rect 270458 220170 300998 220226
rect 301054 220170 301122 220226
rect 301178 220170 331718 220226
rect 331774 220170 331842 220226
rect 331898 220170 362438 220226
rect 362494 220170 362562 220226
rect 362618 220170 393158 220226
rect 393214 220170 393282 220226
rect 393338 220170 423878 220226
rect 423934 220170 424002 220226
rect 424058 220170 454598 220226
rect 454654 220170 454722 220226
rect 454778 220170 485318 220226
rect 485374 220170 485442 220226
rect 485498 220170 516038 220226
rect 516094 220170 516162 220226
rect 516218 220170 525250 220226
rect 525306 220170 525374 220226
rect 525430 220170 525498 220226
rect 525554 220170 525622 220226
rect 525678 220170 543250 220226
rect 543306 220170 543374 220226
rect 543430 220170 543498 220226
rect 543554 220170 543622 220226
rect 543678 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 24518 220102
rect 24574 220046 24642 220102
rect 24698 220046 55238 220102
rect 55294 220046 55362 220102
rect 55418 220046 85958 220102
rect 86014 220046 86082 220102
rect 86138 220046 116678 220102
rect 116734 220046 116802 220102
rect 116858 220046 147398 220102
rect 147454 220046 147522 220102
rect 147578 220046 178118 220102
rect 178174 220046 178242 220102
rect 178298 220046 208838 220102
rect 208894 220046 208962 220102
rect 209018 220046 239558 220102
rect 239614 220046 239682 220102
rect 239738 220046 270278 220102
rect 270334 220046 270402 220102
rect 270458 220046 300998 220102
rect 301054 220046 301122 220102
rect 301178 220046 331718 220102
rect 331774 220046 331842 220102
rect 331898 220046 362438 220102
rect 362494 220046 362562 220102
rect 362618 220046 393158 220102
rect 393214 220046 393282 220102
rect 393338 220046 423878 220102
rect 423934 220046 424002 220102
rect 424058 220046 454598 220102
rect 454654 220046 454722 220102
rect 454778 220046 485318 220102
rect 485374 220046 485442 220102
rect 485498 220046 516038 220102
rect 516094 220046 516162 220102
rect 516218 220046 525250 220102
rect 525306 220046 525374 220102
rect 525430 220046 525498 220102
rect 525554 220046 525622 220102
rect 525678 220046 543250 220102
rect 543306 220046 543374 220102
rect 543430 220046 543498 220102
rect 543554 220046 543622 220102
rect 543678 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 24518 219978
rect 24574 219922 24642 219978
rect 24698 219922 55238 219978
rect 55294 219922 55362 219978
rect 55418 219922 85958 219978
rect 86014 219922 86082 219978
rect 86138 219922 116678 219978
rect 116734 219922 116802 219978
rect 116858 219922 147398 219978
rect 147454 219922 147522 219978
rect 147578 219922 178118 219978
rect 178174 219922 178242 219978
rect 178298 219922 208838 219978
rect 208894 219922 208962 219978
rect 209018 219922 239558 219978
rect 239614 219922 239682 219978
rect 239738 219922 270278 219978
rect 270334 219922 270402 219978
rect 270458 219922 300998 219978
rect 301054 219922 301122 219978
rect 301178 219922 331718 219978
rect 331774 219922 331842 219978
rect 331898 219922 362438 219978
rect 362494 219922 362562 219978
rect 362618 219922 393158 219978
rect 393214 219922 393282 219978
rect 393338 219922 423878 219978
rect 423934 219922 424002 219978
rect 424058 219922 454598 219978
rect 454654 219922 454722 219978
rect 454778 219922 485318 219978
rect 485374 219922 485442 219978
rect 485498 219922 516038 219978
rect 516094 219922 516162 219978
rect 516218 219922 525250 219978
rect 525306 219922 525374 219978
rect 525430 219922 525498 219978
rect 525554 219922 525622 219978
rect 525678 219922 543250 219978
rect 543306 219922 543374 219978
rect 543430 219922 543498 219978
rect 543554 219922 543622 219978
rect 543678 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 39878 208350
rect 39934 208294 40002 208350
rect 40058 208294 70598 208350
rect 70654 208294 70722 208350
rect 70778 208294 101318 208350
rect 101374 208294 101442 208350
rect 101498 208294 132038 208350
rect 132094 208294 132162 208350
rect 132218 208294 162758 208350
rect 162814 208294 162882 208350
rect 162938 208294 193478 208350
rect 193534 208294 193602 208350
rect 193658 208294 224198 208350
rect 224254 208294 224322 208350
rect 224378 208294 254918 208350
rect 254974 208294 255042 208350
rect 255098 208294 285638 208350
rect 285694 208294 285762 208350
rect 285818 208294 316358 208350
rect 316414 208294 316482 208350
rect 316538 208294 347078 208350
rect 347134 208294 347202 208350
rect 347258 208294 377798 208350
rect 377854 208294 377922 208350
rect 377978 208294 408518 208350
rect 408574 208294 408642 208350
rect 408698 208294 439238 208350
rect 439294 208294 439362 208350
rect 439418 208294 469958 208350
rect 470014 208294 470082 208350
rect 470138 208294 500678 208350
rect 500734 208294 500802 208350
rect 500858 208294 528970 208350
rect 529026 208294 529094 208350
rect 529150 208294 529218 208350
rect 529274 208294 529342 208350
rect 529398 208294 546970 208350
rect 547026 208294 547094 208350
rect 547150 208294 547218 208350
rect 547274 208294 547342 208350
rect 547398 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 39878 208226
rect 39934 208170 40002 208226
rect 40058 208170 70598 208226
rect 70654 208170 70722 208226
rect 70778 208170 101318 208226
rect 101374 208170 101442 208226
rect 101498 208170 132038 208226
rect 132094 208170 132162 208226
rect 132218 208170 162758 208226
rect 162814 208170 162882 208226
rect 162938 208170 193478 208226
rect 193534 208170 193602 208226
rect 193658 208170 224198 208226
rect 224254 208170 224322 208226
rect 224378 208170 254918 208226
rect 254974 208170 255042 208226
rect 255098 208170 285638 208226
rect 285694 208170 285762 208226
rect 285818 208170 316358 208226
rect 316414 208170 316482 208226
rect 316538 208170 347078 208226
rect 347134 208170 347202 208226
rect 347258 208170 377798 208226
rect 377854 208170 377922 208226
rect 377978 208170 408518 208226
rect 408574 208170 408642 208226
rect 408698 208170 439238 208226
rect 439294 208170 439362 208226
rect 439418 208170 469958 208226
rect 470014 208170 470082 208226
rect 470138 208170 500678 208226
rect 500734 208170 500802 208226
rect 500858 208170 528970 208226
rect 529026 208170 529094 208226
rect 529150 208170 529218 208226
rect 529274 208170 529342 208226
rect 529398 208170 546970 208226
rect 547026 208170 547094 208226
rect 547150 208170 547218 208226
rect 547274 208170 547342 208226
rect 547398 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 39878 208102
rect 39934 208046 40002 208102
rect 40058 208046 70598 208102
rect 70654 208046 70722 208102
rect 70778 208046 101318 208102
rect 101374 208046 101442 208102
rect 101498 208046 132038 208102
rect 132094 208046 132162 208102
rect 132218 208046 162758 208102
rect 162814 208046 162882 208102
rect 162938 208046 193478 208102
rect 193534 208046 193602 208102
rect 193658 208046 224198 208102
rect 224254 208046 224322 208102
rect 224378 208046 254918 208102
rect 254974 208046 255042 208102
rect 255098 208046 285638 208102
rect 285694 208046 285762 208102
rect 285818 208046 316358 208102
rect 316414 208046 316482 208102
rect 316538 208046 347078 208102
rect 347134 208046 347202 208102
rect 347258 208046 377798 208102
rect 377854 208046 377922 208102
rect 377978 208046 408518 208102
rect 408574 208046 408642 208102
rect 408698 208046 439238 208102
rect 439294 208046 439362 208102
rect 439418 208046 469958 208102
rect 470014 208046 470082 208102
rect 470138 208046 500678 208102
rect 500734 208046 500802 208102
rect 500858 208046 528970 208102
rect 529026 208046 529094 208102
rect 529150 208046 529218 208102
rect 529274 208046 529342 208102
rect 529398 208046 546970 208102
rect 547026 208046 547094 208102
rect 547150 208046 547218 208102
rect 547274 208046 547342 208102
rect 547398 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 39878 207978
rect 39934 207922 40002 207978
rect 40058 207922 70598 207978
rect 70654 207922 70722 207978
rect 70778 207922 101318 207978
rect 101374 207922 101442 207978
rect 101498 207922 132038 207978
rect 132094 207922 132162 207978
rect 132218 207922 162758 207978
rect 162814 207922 162882 207978
rect 162938 207922 193478 207978
rect 193534 207922 193602 207978
rect 193658 207922 224198 207978
rect 224254 207922 224322 207978
rect 224378 207922 254918 207978
rect 254974 207922 255042 207978
rect 255098 207922 285638 207978
rect 285694 207922 285762 207978
rect 285818 207922 316358 207978
rect 316414 207922 316482 207978
rect 316538 207922 347078 207978
rect 347134 207922 347202 207978
rect 347258 207922 377798 207978
rect 377854 207922 377922 207978
rect 377978 207922 408518 207978
rect 408574 207922 408642 207978
rect 408698 207922 439238 207978
rect 439294 207922 439362 207978
rect 439418 207922 469958 207978
rect 470014 207922 470082 207978
rect 470138 207922 500678 207978
rect 500734 207922 500802 207978
rect 500858 207922 528970 207978
rect 529026 207922 529094 207978
rect 529150 207922 529218 207978
rect 529274 207922 529342 207978
rect 529398 207922 546970 207978
rect 547026 207922 547094 207978
rect 547150 207922 547218 207978
rect 547274 207922 547342 207978
rect 547398 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 24518 202350
rect 24574 202294 24642 202350
rect 24698 202294 55238 202350
rect 55294 202294 55362 202350
rect 55418 202294 85958 202350
rect 86014 202294 86082 202350
rect 86138 202294 116678 202350
rect 116734 202294 116802 202350
rect 116858 202294 147398 202350
rect 147454 202294 147522 202350
rect 147578 202294 178118 202350
rect 178174 202294 178242 202350
rect 178298 202294 208838 202350
rect 208894 202294 208962 202350
rect 209018 202294 239558 202350
rect 239614 202294 239682 202350
rect 239738 202294 270278 202350
rect 270334 202294 270402 202350
rect 270458 202294 300998 202350
rect 301054 202294 301122 202350
rect 301178 202294 331718 202350
rect 331774 202294 331842 202350
rect 331898 202294 362438 202350
rect 362494 202294 362562 202350
rect 362618 202294 393158 202350
rect 393214 202294 393282 202350
rect 393338 202294 423878 202350
rect 423934 202294 424002 202350
rect 424058 202294 454598 202350
rect 454654 202294 454722 202350
rect 454778 202294 485318 202350
rect 485374 202294 485442 202350
rect 485498 202294 516038 202350
rect 516094 202294 516162 202350
rect 516218 202294 525250 202350
rect 525306 202294 525374 202350
rect 525430 202294 525498 202350
rect 525554 202294 525622 202350
rect 525678 202294 543250 202350
rect 543306 202294 543374 202350
rect 543430 202294 543498 202350
rect 543554 202294 543622 202350
rect 543678 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 24518 202226
rect 24574 202170 24642 202226
rect 24698 202170 55238 202226
rect 55294 202170 55362 202226
rect 55418 202170 85958 202226
rect 86014 202170 86082 202226
rect 86138 202170 116678 202226
rect 116734 202170 116802 202226
rect 116858 202170 147398 202226
rect 147454 202170 147522 202226
rect 147578 202170 178118 202226
rect 178174 202170 178242 202226
rect 178298 202170 208838 202226
rect 208894 202170 208962 202226
rect 209018 202170 239558 202226
rect 239614 202170 239682 202226
rect 239738 202170 270278 202226
rect 270334 202170 270402 202226
rect 270458 202170 300998 202226
rect 301054 202170 301122 202226
rect 301178 202170 331718 202226
rect 331774 202170 331842 202226
rect 331898 202170 362438 202226
rect 362494 202170 362562 202226
rect 362618 202170 393158 202226
rect 393214 202170 393282 202226
rect 393338 202170 423878 202226
rect 423934 202170 424002 202226
rect 424058 202170 454598 202226
rect 454654 202170 454722 202226
rect 454778 202170 485318 202226
rect 485374 202170 485442 202226
rect 485498 202170 516038 202226
rect 516094 202170 516162 202226
rect 516218 202170 525250 202226
rect 525306 202170 525374 202226
rect 525430 202170 525498 202226
rect 525554 202170 525622 202226
rect 525678 202170 543250 202226
rect 543306 202170 543374 202226
rect 543430 202170 543498 202226
rect 543554 202170 543622 202226
rect 543678 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 24518 202102
rect 24574 202046 24642 202102
rect 24698 202046 55238 202102
rect 55294 202046 55362 202102
rect 55418 202046 85958 202102
rect 86014 202046 86082 202102
rect 86138 202046 116678 202102
rect 116734 202046 116802 202102
rect 116858 202046 147398 202102
rect 147454 202046 147522 202102
rect 147578 202046 178118 202102
rect 178174 202046 178242 202102
rect 178298 202046 208838 202102
rect 208894 202046 208962 202102
rect 209018 202046 239558 202102
rect 239614 202046 239682 202102
rect 239738 202046 270278 202102
rect 270334 202046 270402 202102
rect 270458 202046 300998 202102
rect 301054 202046 301122 202102
rect 301178 202046 331718 202102
rect 331774 202046 331842 202102
rect 331898 202046 362438 202102
rect 362494 202046 362562 202102
rect 362618 202046 393158 202102
rect 393214 202046 393282 202102
rect 393338 202046 423878 202102
rect 423934 202046 424002 202102
rect 424058 202046 454598 202102
rect 454654 202046 454722 202102
rect 454778 202046 485318 202102
rect 485374 202046 485442 202102
rect 485498 202046 516038 202102
rect 516094 202046 516162 202102
rect 516218 202046 525250 202102
rect 525306 202046 525374 202102
rect 525430 202046 525498 202102
rect 525554 202046 525622 202102
rect 525678 202046 543250 202102
rect 543306 202046 543374 202102
rect 543430 202046 543498 202102
rect 543554 202046 543622 202102
rect 543678 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 24518 201978
rect 24574 201922 24642 201978
rect 24698 201922 55238 201978
rect 55294 201922 55362 201978
rect 55418 201922 85958 201978
rect 86014 201922 86082 201978
rect 86138 201922 116678 201978
rect 116734 201922 116802 201978
rect 116858 201922 147398 201978
rect 147454 201922 147522 201978
rect 147578 201922 178118 201978
rect 178174 201922 178242 201978
rect 178298 201922 208838 201978
rect 208894 201922 208962 201978
rect 209018 201922 239558 201978
rect 239614 201922 239682 201978
rect 239738 201922 270278 201978
rect 270334 201922 270402 201978
rect 270458 201922 300998 201978
rect 301054 201922 301122 201978
rect 301178 201922 331718 201978
rect 331774 201922 331842 201978
rect 331898 201922 362438 201978
rect 362494 201922 362562 201978
rect 362618 201922 393158 201978
rect 393214 201922 393282 201978
rect 393338 201922 423878 201978
rect 423934 201922 424002 201978
rect 424058 201922 454598 201978
rect 454654 201922 454722 201978
rect 454778 201922 485318 201978
rect 485374 201922 485442 201978
rect 485498 201922 516038 201978
rect 516094 201922 516162 201978
rect 516218 201922 525250 201978
rect 525306 201922 525374 201978
rect 525430 201922 525498 201978
rect 525554 201922 525622 201978
rect 525678 201922 543250 201978
rect 543306 201922 543374 201978
rect 543430 201922 543498 201978
rect 543554 201922 543622 201978
rect 543678 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 39878 190350
rect 39934 190294 40002 190350
rect 40058 190294 70598 190350
rect 70654 190294 70722 190350
rect 70778 190294 101318 190350
rect 101374 190294 101442 190350
rect 101498 190294 132038 190350
rect 132094 190294 132162 190350
rect 132218 190294 162758 190350
rect 162814 190294 162882 190350
rect 162938 190294 193478 190350
rect 193534 190294 193602 190350
rect 193658 190294 224198 190350
rect 224254 190294 224322 190350
rect 224378 190294 254918 190350
rect 254974 190294 255042 190350
rect 255098 190294 285638 190350
rect 285694 190294 285762 190350
rect 285818 190294 316358 190350
rect 316414 190294 316482 190350
rect 316538 190294 347078 190350
rect 347134 190294 347202 190350
rect 347258 190294 377798 190350
rect 377854 190294 377922 190350
rect 377978 190294 408518 190350
rect 408574 190294 408642 190350
rect 408698 190294 439238 190350
rect 439294 190294 439362 190350
rect 439418 190294 469958 190350
rect 470014 190294 470082 190350
rect 470138 190294 500678 190350
rect 500734 190294 500802 190350
rect 500858 190294 528970 190350
rect 529026 190294 529094 190350
rect 529150 190294 529218 190350
rect 529274 190294 529342 190350
rect 529398 190294 546970 190350
rect 547026 190294 547094 190350
rect 547150 190294 547218 190350
rect 547274 190294 547342 190350
rect 547398 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 39878 190226
rect 39934 190170 40002 190226
rect 40058 190170 70598 190226
rect 70654 190170 70722 190226
rect 70778 190170 101318 190226
rect 101374 190170 101442 190226
rect 101498 190170 132038 190226
rect 132094 190170 132162 190226
rect 132218 190170 162758 190226
rect 162814 190170 162882 190226
rect 162938 190170 193478 190226
rect 193534 190170 193602 190226
rect 193658 190170 224198 190226
rect 224254 190170 224322 190226
rect 224378 190170 254918 190226
rect 254974 190170 255042 190226
rect 255098 190170 285638 190226
rect 285694 190170 285762 190226
rect 285818 190170 316358 190226
rect 316414 190170 316482 190226
rect 316538 190170 347078 190226
rect 347134 190170 347202 190226
rect 347258 190170 377798 190226
rect 377854 190170 377922 190226
rect 377978 190170 408518 190226
rect 408574 190170 408642 190226
rect 408698 190170 439238 190226
rect 439294 190170 439362 190226
rect 439418 190170 469958 190226
rect 470014 190170 470082 190226
rect 470138 190170 500678 190226
rect 500734 190170 500802 190226
rect 500858 190170 528970 190226
rect 529026 190170 529094 190226
rect 529150 190170 529218 190226
rect 529274 190170 529342 190226
rect 529398 190170 546970 190226
rect 547026 190170 547094 190226
rect 547150 190170 547218 190226
rect 547274 190170 547342 190226
rect 547398 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 39878 190102
rect 39934 190046 40002 190102
rect 40058 190046 70598 190102
rect 70654 190046 70722 190102
rect 70778 190046 101318 190102
rect 101374 190046 101442 190102
rect 101498 190046 132038 190102
rect 132094 190046 132162 190102
rect 132218 190046 162758 190102
rect 162814 190046 162882 190102
rect 162938 190046 193478 190102
rect 193534 190046 193602 190102
rect 193658 190046 224198 190102
rect 224254 190046 224322 190102
rect 224378 190046 254918 190102
rect 254974 190046 255042 190102
rect 255098 190046 285638 190102
rect 285694 190046 285762 190102
rect 285818 190046 316358 190102
rect 316414 190046 316482 190102
rect 316538 190046 347078 190102
rect 347134 190046 347202 190102
rect 347258 190046 377798 190102
rect 377854 190046 377922 190102
rect 377978 190046 408518 190102
rect 408574 190046 408642 190102
rect 408698 190046 439238 190102
rect 439294 190046 439362 190102
rect 439418 190046 469958 190102
rect 470014 190046 470082 190102
rect 470138 190046 500678 190102
rect 500734 190046 500802 190102
rect 500858 190046 528970 190102
rect 529026 190046 529094 190102
rect 529150 190046 529218 190102
rect 529274 190046 529342 190102
rect 529398 190046 546970 190102
rect 547026 190046 547094 190102
rect 547150 190046 547218 190102
rect 547274 190046 547342 190102
rect 547398 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 39878 189978
rect 39934 189922 40002 189978
rect 40058 189922 70598 189978
rect 70654 189922 70722 189978
rect 70778 189922 101318 189978
rect 101374 189922 101442 189978
rect 101498 189922 132038 189978
rect 132094 189922 132162 189978
rect 132218 189922 162758 189978
rect 162814 189922 162882 189978
rect 162938 189922 193478 189978
rect 193534 189922 193602 189978
rect 193658 189922 224198 189978
rect 224254 189922 224322 189978
rect 224378 189922 254918 189978
rect 254974 189922 255042 189978
rect 255098 189922 285638 189978
rect 285694 189922 285762 189978
rect 285818 189922 316358 189978
rect 316414 189922 316482 189978
rect 316538 189922 347078 189978
rect 347134 189922 347202 189978
rect 347258 189922 377798 189978
rect 377854 189922 377922 189978
rect 377978 189922 408518 189978
rect 408574 189922 408642 189978
rect 408698 189922 439238 189978
rect 439294 189922 439362 189978
rect 439418 189922 469958 189978
rect 470014 189922 470082 189978
rect 470138 189922 500678 189978
rect 500734 189922 500802 189978
rect 500858 189922 528970 189978
rect 529026 189922 529094 189978
rect 529150 189922 529218 189978
rect 529274 189922 529342 189978
rect 529398 189922 546970 189978
rect 547026 189922 547094 189978
rect 547150 189922 547218 189978
rect 547274 189922 547342 189978
rect 547398 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 24518 184350
rect 24574 184294 24642 184350
rect 24698 184294 55238 184350
rect 55294 184294 55362 184350
rect 55418 184294 85958 184350
rect 86014 184294 86082 184350
rect 86138 184294 116678 184350
rect 116734 184294 116802 184350
rect 116858 184294 147398 184350
rect 147454 184294 147522 184350
rect 147578 184294 178118 184350
rect 178174 184294 178242 184350
rect 178298 184294 208838 184350
rect 208894 184294 208962 184350
rect 209018 184294 239558 184350
rect 239614 184294 239682 184350
rect 239738 184294 270278 184350
rect 270334 184294 270402 184350
rect 270458 184294 300998 184350
rect 301054 184294 301122 184350
rect 301178 184294 331718 184350
rect 331774 184294 331842 184350
rect 331898 184294 362438 184350
rect 362494 184294 362562 184350
rect 362618 184294 393158 184350
rect 393214 184294 393282 184350
rect 393338 184294 423878 184350
rect 423934 184294 424002 184350
rect 424058 184294 454598 184350
rect 454654 184294 454722 184350
rect 454778 184294 485318 184350
rect 485374 184294 485442 184350
rect 485498 184294 516038 184350
rect 516094 184294 516162 184350
rect 516218 184294 525250 184350
rect 525306 184294 525374 184350
rect 525430 184294 525498 184350
rect 525554 184294 525622 184350
rect 525678 184294 543250 184350
rect 543306 184294 543374 184350
rect 543430 184294 543498 184350
rect 543554 184294 543622 184350
rect 543678 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 24518 184226
rect 24574 184170 24642 184226
rect 24698 184170 55238 184226
rect 55294 184170 55362 184226
rect 55418 184170 85958 184226
rect 86014 184170 86082 184226
rect 86138 184170 116678 184226
rect 116734 184170 116802 184226
rect 116858 184170 147398 184226
rect 147454 184170 147522 184226
rect 147578 184170 178118 184226
rect 178174 184170 178242 184226
rect 178298 184170 208838 184226
rect 208894 184170 208962 184226
rect 209018 184170 239558 184226
rect 239614 184170 239682 184226
rect 239738 184170 270278 184226
rect 270334 184170 270402 184226
rect 270458 184170 300998 184226
rect 301054 184170 301122 184226
rect 301178 184170 331718 184226
rect 331774 184170 331842 184226
rect 331898 184170 362438 184226
rect 362494 184170 362562 184226
rect 362618 184170 393158 184226
rect 393214 184170 393282 184226
rect 393338 184170 423878 184226
rect 423934 184170 424002 184226
rect 424058 184170 454598 184226
rect 454654 184170 454722 184226
rect 454778 184170 485318 184226
rect 485374 184170 485442 184226
rect 485498 184170 516038 184226
rect 516094 184170 516162 184226
rect 516218 184170 525250 184226
rect 525306 184170 525374 184226
rect 525430 184170 525498 184226
rect 525554 184170 525622 184226
rect 525678 184170 543250 184226
rect 543306 184170 543374 184226
rect 543430 184170 543498 184226
rect 543554 184170 543622 184226
rect 543678 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 24518 184102
rect 24574 184046 24642 184102
rect 24698 184046 55238 184102
rect 55294 184046 55362 184102
rect 55418 184046 85958 184102
rect 86014 184046 86082 184102
rect 86138 184046 116678 184102
rect 116734 184046 116802 184102
rect 116858 184046 147398 184102
rect 147454 184046 147522 184102
rect 147578 184046 178118 184102
rect 178174 184046 178242 184102
rect 178298 184046 208838 184102
rect 208894 184046 208962 184102
rect 209018 184046 239558 184102
rect 239614 184046 239682 184102
rect 239738 184046 270278 184102
rect 270334 184046 270402 184102
rect 270458 184046 300998 184102
rect 301054 184046 301122 184102
rect 301178 184046 331718 184102
rect 331774 184046 331842 184102
rect 331898 184046 362438 184102
rect 362494 184046 362562 184102
rect 362618 184046 393158 184102
rect 393214 184046 393282 184102
rect 393338 184046 423878 184102
rect 423934 184046 424002 184102
rect 424058 184046 454598 184102
rect 454654 184046 454722 184102
rect 454778 184046 485318 184102
rect 485374 184046 485442 184102
rect 485498 184046 516038 184102
rect 516094 184046 516162 184102
rect 516218 184046 525250 184102
rect 525306 184046 525374 184102
rect 525430 184046 525498 184102
rect 525554 184046 525622 184102
rect 525678 184046 543250 184102
rect 543306 184046 543374 184102
rect 543430 184046 543498 184102
rect 543554 184046 543622 184102
rect 543678 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 24518 183978
rect 24574 183922 24642 183978
rect 24698 183922 55238 183978
rect 55294 183922 55362 183978
rect 55418 183922 85958 183978
rect 86014 183922 86082 183978
rect 86138 183922 116678 183978
rect 116734 183922 116802 183978
rect 116858 183922 147398 183978
rect 147454 183922 147522 183978
rect 147578 183922 178118 183978
rect 178174 183922 178242 183978
rect 178298 183922 208838 183978
rect 208894 183922 208962 183978
rect 209018 183922 239558 183978
rect 239614 183922 239682 183978
rect 239738 183922 270278 183978
rect 270334 183922 270402 183978
rect 270458 183922 300998 183978
rect 301054 183922 301122 183978
rect 301178 183922 331718 183978
rect 331774 183922 331842 183978
rect 331898 183922 362438 183978
rect 362494 183922 362562 183978
rect 362618 183922 393158 183978
rect 393214 183922 393282 183978
rect 393338 183922 423878 183978
rect 423934 183922 424002 183978
rect 424058 183922 454598 183978
rect 454654 183922 454722 183978
rect 454778 183922 485318 183978
rect 485374 183922 485442 183978
rect 485498 183922 516038 183978
rect 516094 183922 516162 183978
rect 516218 183922 525250 183978
rect 525306 183922 525374 183978
rect 525430 183922 525498 183978
rect 525554 183922 525622 183978
rect 525678 183922 543250 183978
rect 543306 183922 543374 183978
rect 543430 183922 543498 183978
rect 543554 183922 543622 183978
rect 543678 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 39878 172350
rect 39934 172294 40002 172350
rect 40058 172294 70598 172350
rect 70654 172294 70722 172350
rect 70778 172294 101318 172350
rect 101374 172294 101442 172350
rect 101498 172294 132038 172350
rect 132094 172294 132162 172350
rect 132218 172294 162758 172350
rect 162814 172294 162882 172350
rect 162938 172294 193478 172350
rect 193534 172294 193602 172350
rect 193658 172294 224198 172350
rect 224254 172294 224322 172350
rect 224378 172294 254918 172350
rect 254974 172294 255042 172350
rect 255098 172294 285638 172350
rect 285694 172294 285762 172350
rect 285818 172294 316358 172350
rect 316414 172294 316482 172350
rect 316538 172294 347078 172350
rect 347134 172294 347202 172350
rect 347258 172294 377798 172350
rect 377854 172294 377922 172350
rect 377978 172294 408518 172350
rect 408574 172294 408642 172350
rect 408698 172294 439238 172350
rect 439294 172294 439362 172350
rect 439418 172294 469958 172350
rect 470014 172294 470082 172350
rect 470138 172294 500678 172350
rect 500734 172294 500802 172350
rect 500858 172294 528970 172350
rect 529026 172294 529094 172350
rect 529150 172294 529218 172350
rect 529274 172294 529342 172350
rect 529398 172294 546970 172350
rect 547026 172294 547094 172350
rect 547150 172294 547218 172350
rect 547274 172294 547342 172350
rect 547398 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 39878 172226
rect 39934 172170 40002 172226
rect 40058 172170 70598 172226
rect 70654 172170 70722 172226
rect 70778 172170 101318 172226
rect 101374 172170 101442 172226
rect 101498 172170 132038 172226
rect 132094 172170 132162 172226
rect 132218 172170 162758 172226
rect 162814 172170 162882 172226
rect 162938 172170 193478 172226
rect 193534 172170 193602 172226
rect 193658 172170 224198 172226
rect 224254 172170 224322 172226
rect 224378 172170 254918 172226
rect 254974 172170 255042 172226
rect 255098 172170 285638 172226
rect 285694 172170 285762 172226
rect 285818 172170 316358 172226
rect 316414 172170 316482 172226
rect 316538 172170 347078 172226
rect 347134 172170 347202 172226
rect 347258 172170 377798 172226
rect 377854 172170 377922 172226
rect 377978 172170 408518 172226
rect 408574 172170 408642 172226
rect 408698 172170 439238 172226
rect 439294 172170 439362 172226
rect 439418 172170 469958 172226
rect 470014 172170 470082 172226
rect 470138 172170 500678 172226
rect 500734 172170 500802 172226
rect 500858 172170 528970 172226
rect 529026 172170 529094 172226
rect 529150 172170 529218 172226
rect 529274 172170 529342 172226
rect 529398 172170 546970 172226
rect 547026 172170 547094 172226
rect 547150 172170 547218 172226
rect 547274 172170 547342 172226
rect 547398 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 39878 172102
rect 39934 172046 40002 172102
rect 40058 172046 70598 172102
rect 70654 172046 70722 172102
rect 70778 172046 101318 172102
rect 101374 172046 101442 172102
rect 101498 172046 132038 172102
rect 132094 172046 132162 172102
rect 132218 172046 162758 172102
rect 162814 172046 162882 172102
rect 162938 172046 193478 172102
rect 193534 172046 193602 172102
rect 193658 172046 224198 172102
rect 224254 172046 224322 172102
rect 224378 172046 254918 172102
rect 254974 172046 255042 172102
rect 255098 172046 285638 172102
rect 285694 172046 285762 172102
rect 285818 172046 316358 172102
rect 316414 172046 316482 172102
rect 316538 172046 347078 172102
rect 347134 172046 347202 172102
rect 347258 172046 377798 172102
rect 377854 172046 377922 172102
rect 377978 172046 408518 172102
rect 408574 172046 408642 172102
rect 408698 172046 439238 172102
rect 439294 172046 439362 172102
rect 439418 172046 469958 172102
rect 470014 172046 470082 172102
rect 470138 172046 500678 172102
rect 500734 172046 500802 172102
rect 500858 172046 528970 172102
rect 529026 172046 529094 172102
rect 529150 172046 529218 172102
rect 529274 172046 529342 172102
rect 529398 172046 546970 172102
rect 547026 172046 547094 172102
rect 547150 172046 547218 172102
rect 547274 172046 547342 172102
rect 547398 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 39878 171978
rect 39934 171922 40002 171978
rect 40058 171922 70598 171978
rect 70654 171922 70722 171978
rect 70778 171922 101318 171978
rect 101374 171922 101442 171978
rect 101498 171922 132038 171978
rect 132094 171922 132162 171978
rect 132218 171922 162758 171978
rect 162814 171922 162882 171978
rect 162938 171922 193478 171978
rect 193534 171922 193602 171978
rect 193658 171922 224198 171978
rect 224254 171922 224322 171978
rect 224378 171922 254918 171978
rect 254974 171922 255042 171978
rect 255098 171922 285638 171978
rect 285694 171922 285762 171978
rect 285818 171922 316358 171978
rect 316414 171922 316482 171978
rect 316538 171922 347078 171978
rect 347134 171922 347202 171978
rect 347258 171922 377798 171978
rect 377854 171922 377922 171978
rect 377978 171922 408518 171978
rect 408574 171922 408642 171978
rect 408698 171922 439238 171978
rect 439294 171922 439362 171978
rect 439418 171922 469958 171978
rect 470014 171922 470082 171978
rect 470138 171922 500678 171978
rect 500734 171922 500802 171978
rect 500858 171922 528970 171978
rect 529026 171922 529094 171978
rect 529150 171922 529218 171978
rect 529274 171922 529342 171978
rect 529398 171922 546970 171978
rect 547026 171922 547094 171978
rect 547150 171922 547218 171978
rect 547274 171922 547342 171978
rect 547398 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 24518 166350
rect 24574 166294 24642 166350
rect 24698 166294 55238 166350
rect 55294 166294 55362 166350
rect 55418 166294 85958 166350
rect 86014 166294 86082 166350
rect 86138 166294 116678 166350
rect 116734 166294 116802 166350
rect 116858 166294 147398 166350
rect 147454 166294 147522 166350
rect 147578 166294 178118 166350
rect 178174 166294 178242 166350
rect 178298 166294 208838 166350
rect 208894 166294 208962 166350
rect 209018 166294 239558 166350
rect 239614 166294 239682 166350
rect 239738 166294 270278 166350
rect 270334 166294 270402 166350
rect 270458 166294 300998 166350
rect 301054 166294 301122 166350
rect 301178 166294 331718 166350
rect 331774 166294 331842 166350
rect 331898 166294 362438 166350
rect 362494 166294 362562 166350
rect 362618 166294 393158 166350
rect 393214 166294 393282 166350
rect 393338 166294 423878 166350
rect 423934 166294 424002 166350
rect 424058 166294 454598 166350
rect 454654 166294 454722 166350
rect 454778 166294 485318 166350
rect 485374 166294 485442 166350
rect 485498 166294 516038 166350
rect 516094 166294 516162 166350
rect 516218 166294 525250 166350
rect 525306 166294 525374 166350
rect 525430 166294 525498 166350
rect 525554 166294 525622 166350
rect 525678 166294 543250 166350
rect 543306 166294 543374 166350
rect 543430 166294 543498 166350
rect 543554 166294 543622 166350
rect 543678 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 24518 166226
rect 24574 166170 24642 166226
rect 24698 166170 55238 166226
rect 55294 166170 55362 166226
rect 55418 166170 85958 166226
rect 86014 166170 86082 166226
rect 86138 166170 116678 166226
rect 116734 166170 116802 166226
rect 116858 166170 147398 166226
rect 147454 166170 147522 166226
rect 147578 166170 178118 166226
rect 178174 166170 178242 166226
rect 178298 166170 208838 166226
rect 208894 166170 208962 166226
rect 209018 166170 239558 166226
rect 239614 166170 239682 166226
rect 239738 166170 270278 166226
rect 270334 166170 270402 166226
rect 270458 166170 300998 166226
rect 301054 166170 301122 166226
rect 301178 166170 331718 166226
rect 331774 166170 331842 166226
rect 331898 166170 362438 166226
rect 362494 166170 362562 166226
rect 362618 166170 393158 166226
rect 393214 166170 393282 166226
rect 393338 166170 423878 166226
rect 423934 166170 424002 166226
rect 424058 166170 454598 166226
rect 454654 166170 454722 166226
rect 454778 166170 485318 166226
rect 485374 166170 485442 166226
rect 485498 166170 516038 166226
rect 516094 166170 516162 166226
rect 516218 166170 525250 166226
rect 525306 166170 525374 166226
rect 525430 166170 525498 166226
rect 525554 166170 525622 166226
rect 525678 166170 543250 166226
rect 543306 166170 543374 166226
rect 543430 166170 543498 166226
rect 543554 166170 543622 166226
rect 543678 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 24518 166102
rect 24574 166046 24642 166102
rect 24698 166046 55238 166102
rect 55294 166046 55362 166102
rect 55418 166046 85958 166102
rect 86014 166046 86082 166102
rect 86138 166046 116678 166102
rect 116734 166046 116802 166102
rect 116858 166046 147398 166102
rect 147454 166046 147522 166102
rect 147578 166046 178118 166102
rect 178174 166046 178242 166102
rect 178298 166046 208838 166102
rect 208894 166046 208962 166102
rect 209018 166046 239558 166102
rect 239614 166046 239682 166102
rect 239738 166046 270278 166102
rect 270334 166046 270402 166102
rect 270458 166046 300998 166102
rect 301054 166046 301122 166102
rect 301178 166046 331718 166102
rect 331774 166046 331842 166102
rect 331898 166046 362438 166102
rect 362494 166046 362562 166102
rect 362618 166046 393158 166102
rect 393214 166046 393282 166102
rect 393338 166046 423878 166102
rect 423934 166046 424002 166102
rect 424058 166046 454598 166102
rect 454654 166046 454722 166102
rect 454778 166046 485318 166102
rect 485374 166046 485442 166102
rect 485498 166046 516038 166102
rect 516094 166046 516162 166102
rect 516218 166046 525250 166102
rect 525306 166046 525374 166102
rect 525430 166046 525498 166102
rect 525554 166046 525622 166102
rect 525678 166046 543250 166102
rect 543306 166046 543374 166102
rect 543430 166046 543498 166102
rect 543554 166046 543622 166102
rect 543678 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 24518 165978
rect 24574 165922 24642 165978
rect 24698 165922 55238 165978
rect 55294 165922 55362 165978
rect 55418 165922 85958 165978
rect 86014 165922 86082 165978
rect 86138 165922 116678 165978
rect 116734 165922 116802 165978
rect 116858 165922 147398 165978
rect 147454 165922 147522 165978
rect 147578 165922 178118 165978
rect 178174 165922 178242 165978
rect 178298 165922 208838 165978
rect 208894 165922 208962 165978
rect 209018 165922 239558 165978
rect 239614 165922 239682 165978
rect 239738 165922 270278 165978
rect 270334 165922 270402 165978
rect 270458 165922 300998 165978
rect 301054 165922 301122 165978
rect 301178 165922 331718 165978
rect 331774 165922 331842 165978
rect 331898 165922 362438 165978
rect 362494 165922 362562 165978
rect 362618 165922 393158 165978
rect 393214 165922 393282 165978
rect 393338 165922 423878 165978
rect 423934 165922 424002 165978
rect 424058 165922 454598 165978
rect 454654 165922 454722 165978
rect 454778 165922 485318 165978
rect 485374 165922 485442 165978
rect 485498 165922 516038 165978
rect 516094 165922 516162 165978
rect 516218 165922 525250 165978
rect 525306 165922 525374 165978
rect 525430 165922 525498 165978
rect 525554 165922 525622 165978
rect 525678 165922 543250 165978
rect 543306 165922 543374 165978
rect 543430 165922 543498 165978
rect 543554 165922 543622 165978
rect 543678 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 39878 154350
rect 39934 154294 40002 154350
rect 40058 154294 70598 154350
rect 70654 154294 70722 154350
rect 70778 154294 101318 154350
rect 101374 154294 101442 154350
rect 101498 154294 132038 154350
rect 132094 154294 132162 154350
rect 132218 154294 162758 154350
rect 162814 154294 162882 154350
rect 162938 154294 193478 154350
rect 193534 154294 193602 154350
rect 193658 154294 224198 154350
rect 224254 154294 224322 154350
rect 224378 154294 254918 154350
rect 254974 154294 255042 154350
rect 255098 154294 285638 154350
rect 285694 154294 285762 154350
rect 285818 154294 316358 154350
rect 316414 154294 316482 154350
rect 316538 154294 347078 154350
rect 347134 154294 347202 154350
rect 347258 154294 377798 154350
rect 377854 154294 377922 154350
rect 377978 154294 408518 154350
rect 408574 154294 408642 154350
rect 408698 154294 439238 154350
rect 439294 154294 439362 154350
rect 439418 154294 469958 154350
rect 470014 154294 470082 154350
rect 470138 154294 500678 154350
rect 500734 154294 500802 154350
rect 500858 154294 528970 154350
rect 529026 154294 529094 154350
rect 529150 154294 529218 154350
rect 529274 154294 529342 154350
rect 529398 154294 546970 154350
rect 547026 154294 547094 154350
rect 547150 154294 547218 154350
rect 547274 154294 547342 154350
rect 547398 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 39878 154226
rect 39934 154170 40002 154226
rect 40058 154170 70598 154226
rect 70654 154170 70722 154226
rect 70778 154170 101318 154226
rect 101374 154170 101442 154226
rect 101498 154170 132038 154226
rect 132094 154170 132162 154226
rect 132218 154170 162758 154226
rect 162814 154170 162882 154226
rect 162938 154170 193478 154226
rect 193534 154170 193602 154226
rect 193658 154170 224198 154226
rect 224254 154170 224322 154226
rect 224378 154170 254918 154226
rect 254974 154170 255042 154226
rect 255098 154170 285638 154226
rect 285694 154170 285762 154226
rect 285818 154170 316358 154226
rect 316414 154170 316482 154226
rect 316538 154170 347078 154226
rect 347134 154170 347202 154226
rect 347258 154170 377798 154226
rect 377854 154170 377922 154226
rect 377978 154170 408518 154226
rect 408574 154170 408642 154226
rect 408698 154170 439238 154226
rect 439294 154170 439362 154226
rect 439418 154170 469958 154226
rect 470014 154170 470082 154226
rect 470138 154170 500678 154226
rect 500734 154170 500802 154226
rect 500858 154170 528970 154226
rect 529026 154170 529094 154226
rect 529150 154170 529218 154226
rect 529274 154170 529342 154226
rect 529398 154170 546970 154226
rect 547026 154170 547094 154226
rect 547150 154170 547218 154226
rect 547274 154170 547342 154226
rect 547398 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 39878 154102
rect 39934 154046 40002 154102
rect 40058 154046 70598 154102
rect 70654 154046 70722 154102
rect 70778 154046 101318 154102
rect 101374 154046 101442 154102
rect 101498 154046 132038 154102
rect 132094 154046 132162 154102
rect 132218 154046 162758 154102
rect 162814 154046 162882 154102
rect 162938 154046 193478 154102
rect 193534 154046 193602 154102
rect 193658 154046 224198 154102
rect 224254 154046 224322 154102
rect 224378 154046 254918 154102
rect 254974 154046 255042 154102
rect 255098 154046 285638 154102
rect 285694 154046 285762 154102
rect 285818 154046 316358 154102
rect 316414 154046 316482 154102
rect 316538 154046 347078 154102
rect 347134 154046 347202 154102
rect 347258 154046 377798 154102
rect 377854 154046 377922 154102
rect 377978 154046 408518 154102
rect 408574 154046 408642 154102
rect 408698 154046 439238 154102
rect 439294 154046 439362 154102
rect 439418 154046 469958 154102
rect 470014 154046 470082 154102
rect 470138 154046 500678 154102
rect 500734 154046 500802 154102
rect 500858 154046 528970 154102
rect 529026 154046 529094 154102
rect 529150 154046 529218 154102
rect 529274 154046 529342 154102
rect 529398 154046 546970 154102
rect 547026 154046 547094 154102
rect 547150 154046 547218 154102
rect 547274 154046 547342 154102
rect 547398 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 39878 153978
rect 39934 153922 40002 153978
rect 40058 153922 70598 153978
rect 70654 153922 70722 153978
rect 70778 153922 101318 153978
rect 101374 153922 101442 153978
rect 101498 153922 132038 153978
rect 132094 153922 132162 153978
rect 132218 153922 162758 153978
rect 162814 153922 162882 153978
rect 162938 153922 193478 153978
rect 193534 153922 193602 153978
rect 193658 153922 224198 153978
rect 224254 153922 224322 153978
rect 224378 153922 254918 153978
rect 254974 153922 255042 153978
rect 255098 153922 285638 153978
rect 285694 153922 285762 153978
rect 285818 153922 316358 153978
rect 316414 153922 316482 153978
rect 316538 153922 347078 153978
rect 347134 153922 347202 153978
rect 347258 153922 377798 153978
rect 377854 153922 377922 153978
rect 377978 153922 408518 153978
rect 408574 153922 408642 153978
rect 408698 153922 439238 153978
rect 439294 153922 439362 153978
rect 439418 153922 469958 153978
rect 470014 153922 470082 153978
rect 470138 153922 500678 153978
rect 500734 153922 500802 153978
rect 500858 153922 528970 153978
rect 529026 153922 529094 153978
rect 529150 153922 529218 153978
rect 529274 153922 529342 153978
rect 529398 153922 546970 153978
rect 547026 153922 547094 153978
rect 547150 153922 547218 153978
rect 547274 153922 547342 153978
rect 547398 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 24518 148350
rect 24574 148294 24642 148350
rect 24698 148294 55238 148350
rect 55294 148294 55362 148350
rect 55418 148294 85958 148350
rect 86014 148294 86082 148350
rect 86138 148294 116678 148350
rect 116734 148294 116802 148350
rect 116858 148294 147398 148350
rect 147454 148294 147522 148350
rect 147578 148294 178118 148350
rect 178174 148294 178242 148350
rect 178298 148294 208838 148350
rect 208894 148294 208962 148350
rect 209018 148294 239558 148350
rect 239614 148294 239682 148350
rect 239738 148294 270278 148350
rect 270334 148294 270402 148350
rect 270458 148294 300998 148350
rect 301054 148294 301122 148350
rect 301178 148294 331718 148350
rect 331774 148294 331842 148350
rect 331898 148294 362438 148350
rect 362494 148294 362562 148350
rect 362618 148294 393158 148350
rect 393214 148294 393282 148350
rect 393338 148294 423878 148350
rect 423934 148294 424002 148350
rect 424058 148294 454598 148350
rect 454654 148294 454722 148350
rect 454778 148294 485318 148350
rect 485374 148294 485442 148350
rect 485498 148294 516038 148350
rect 516094 148294 516162 148350
rect 516218 148294 525250 148350
rect 525306 148294 525374 148350
rect 525430 148294 525498 148350
rect 525554 148294 525622 148350
rect 525678 148294 543250 148350
rect 543306 148294 543374 148350
rect 543430 148294 543498 148350
rect 543554 148294 543622 148350
rect 543678 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 24518 148226
rect 24574 148170 24642 148226
rect 24698 148170 55238 148226
rect 55294 148170 55362 148226
rect 55418 148170 85958 148226
rect 86014 148170 86082 148226
rect 86138 148170 116678 148226
rect 116734 148170 116802 148226
rect 116858 148170 147398 148226
rect 147454 148170 147522 148226
rect 147578 148170 178118 148226
rect 178174 148170 178242 148226
rect 178298 148170 208838 148226
rect 208894 148170 208962 148226
rect 209018 148170 239558 148226
rect 239614 148170 239682 148226
rect 239738 148170 270278 148226
rect 270334 148170 270402 148226
rect 270458 148170 300998 148226
rect 301054 148170 301122 148226
rect 301178 148170 331718 148226
rect 331774 148170 331842 148226
rect 331898 148170 362438 148226
rect 362494 148170 362562 148226
rect 362618 148170 393158 148226
rect 393214 148170 393282 148226
rect 393338 148170 423878 148226
rect 423934 148170 424002 148226
rect 424058 148170 454598 148226
rect 454654 148170 454722 148226
rect 454778 148170 485318 148226
rect 485374 148170 485442 148226
rect 485498 148170 516038 148226
rect 516094 148170 516162 148226
rect 516218 148170 525250 148226
rect 525306 148170 525374 148226
rect 525430 148170 525498 148226
rect 525554 148170 525622 148226
rect 525678 148170 543250 148226
rect 543306 148170 543374 148226
rect 543430 148170 543498 148226
rect 543554 148170 543622 148226
rect 543678 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 24518 148102
rect 24574 148046 24642 148102
rect 24698 148046 55238 148102
rect 55294 148046 55362 148102
rect 55418 148046 85958 148102
rect 86014 148046 86082 148102
rect 86138 148046 116678 148102
rect 116734 148046 116802 148102
rect 116858 148046 147398 148102
rect 147454 148046 147522 148102
rect 147578 148046 178118 148102
rect 178174 148046 178242 148102
rect 178298 148046 208838 148102
rect 208894 148046 208962 148102
rect 209018 148046 239558 148102
rect 239614 148046 239682 148102
rect 239738 148046 270278 148102
rect 270334 148046 270402 148102
rect 270458 148046 300998 148102
rect 301054 148046 301122 148102
rect 301178 148046 331718 148102
rect 331774 148046 331842 148102
rect 331898 148046 362438 148102
rect 362494 148046 362562 148102
rect 362618 148046 393158 148102
rect 393214 148046 393282 148102
rect 393338 148046 423878 148102
rect 423934 148046 424002 148102
rect 424058 148046 454598 148102
rect 454654 148046 454722 148102
rect 454778 148046 485318 148102
rect 485374 148046 485442 148102
rect 485498 148046 516038 148102
rect 516094 148046 516162 148102
rect 516218 148046 525250 148102
rect 525306 148046 525374 148102
rect 525430 148046 525498 148102
rect 525554 148046 525622 148102
rect 525678 148046 543250 148102
rect 543306 148046 543374 148102
rect 543430 148046 543498 148102
rect 543554 148046 543622 148102
rect 543678 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 24518 147978
rect 24574 147922 24642 147978
rect 24698 147922 55238 147978
rect 55294 147922 55362 147978
rect 55418 147922 85958 147978
rect 86014 147922 86082 147978
rect 86138 147922 116678 147978
rect 116734 147922 116802 147978
rect 116858 147922 147398 147978
rect 147454 147922 147522 147978
rect 147578 147922 178118 147978
rect 178174 147922 178242 147978
rect 178298 147922 208838 147978
rect 208894 147922 208962 147978
rect 209018 147922 239558 147978
rect 239614 147922 239682 147978
rect 239738 147922 270278 147978
rect 270334 147922 270402 147978
rect 270458 147922 300998 147978
rect 301054 147922 301122 147978
rect 301178 147922 331718 147978
rect 331774 147922 331842 147978
rect 331898 147922 362438 147978
rect 362494 147922 362562 147978
rect 362618 147922 393158 147978
rect 393214 147922 393282 147978
rect 393338 147922 423878 147978
rect 423934 147922 424002 147978
rect 424058 147922 454598 147978
rect 454654 147922 454722 147978
rect 454778 147922 485318 147978
rect 485374 147922 485442 147978
rect 485498 147922 516038 147978
rect 516094 147922 516162 147978
rect 516218 147922 525250 147978
rect 525306 147922 525374 147978
rect 525430 147922 525498 147978
rect 525554 147922 525622 147978
rect 525678 147922 543250 147978
rect 543306 147922 543374 147978
rect 543430 147922 543498 147978
rect 543554 147922 543622 147978
rect 543678 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 39878 136350
rect 39934 136294 40002 136350
rect 40058 136294 70598 136350
rect 70654 136294 70722 136350
rect 70778 136294 101318 136350
rect 101374 136294 101442 136350
rect 101498 136294 132038 136350
rect 132094 136294 132162 136350
rect 132218 136294 162758 136350
rect 162814 136294 162882 136350
rect 162938 136294 193478 136350
rect 193534 136294 193602 136350
rect 193658 136294 224198 136350
rect 224254 136294 224322 136350
rect 224378 136294 254918 136350
rect 254974 136294 255042 136350
rect 255098 136294 285638 136350
rect 285694 136294 285762 136350
rect 285818 136294 316358 136350
rect 316414 136294 316482 136350
rect 316538 136294 347078 136350
rect 347134 136294 347202 136350
rect 347258 136294 377798 136350
rect 377854 136294 377922 136350
rect 377978 136294 408518 136350
rect 408574 136294 408642 136350
rect 408698 136294 439238 136350
rect 439294 136294 439362 136350
rect 439418 136294 469958 136350
rect 470014 136294 470082 136350
rect 470138 136294 500678 136350
rect 500734 136294 500802 136350
rect 500858 136294 528970 136350
rect 529026 136294 529094 136350
rect 529150 136294 529218 136350
rect 529274 136294 529342 136350
rect 529398 136294 546970 136350
rect 547026 136294 547094 136350
rect 547150 136294 547218 136350
rect 547274 136294 547342 136350
rect 547398 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 39878 136226
rect 39934 136170 40002 136226
rect 40058 136170 70598 136226
rect 70654 136170 70722 136226
rect 70778 136170 101318 136226
rect 101374 136170 101442 136226
rect 101498 136170 132038 136226
rect 132094 136170 132162 136226
rect 132218 136170 162758 136226
rect 162814 136170 162882 136226
rect 162938 136170 193478 136226
rect 193534 136170 193602 136226
rect 193658 136170 224198 136226
rect 224254 136170 224322 136226
rect 224378 136170 254918 136226
rect 254974 136170 255042 136226
rect 255098 136170 285638 136226
rect 285694 136170 285762 136226
rect 285818 136170 316358 136226
rect 316414 136170 316482 136226
rect 316538 136170 347078 136226
rect 347134 136170 347202 136226
rect 347258 136170 377798 136226
rect 377854 136170 377922 136226
rect 377978 136170 408518 136226
rect 408574 136170 408642 136226
rect 408698 136170 439238 136226
rect 439294 136170 439362 136226
rect 439418 136170 469958 136226
rect 470014 136170 470082 136226
rect 470138 136170 500678 136226
rect 500734 136170 500802 136226
rect 500858 136170 528970 136226
rect 529026 136170 529094 136226
rect 529150 136170 529218 136226
rect 529274 136170 529342 136226
rect 529398 136170 546970 136226
rect 547026 136170 547094 136226
rect 547150 136170 547218 136226
rect 547274 136170 547342 136226
rect 547398 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 39878 136102
rect 39934 136046 40002 136102
rect 40058 136046 70598 136102
rect 70654 136046 70722 136102
rect 70778 136046 101318 136102
rect 101374 136046 101442 136102
rect 101498 136046 132038 136102
rect 132094 136046 132162 136102
rect 132218 136046 162758 136102
rect 162814 136046 162882 136102
rect 162938 136046 193478 136102
rect 193534 136046 193602 136102
rect 193658 136046 224198 136102
rect 224254 136046 224322 136102
rect 224378 136046 254918 136102
rect 254974 136046 255042 136102
rect 255098 136046 285638 136102
rect 285694 136046 285762 136102
rect 285818 136046 316358 136102
rect 316414 136046 316482 136102
rect 316538 136046 347078 136102
rect 347134 136046 347202 136102
rect 347258 136046 377798 136102
rect 377854 136046 377922 136102
rect 377978 136046 408518 136102
rect 408574 136046 408642 136102
rect 408698 136046 439238 136102
rect 439294 136046 439362 136102
rect 439418 136046 469958 136102
rect 470014 136046 470082 136102
rect 470138 136046 500678 136102
rect 500734 136046 500802 136102
rect 500858 136046 528970 136102
rect 529026 136046 529094 136102
rect 529150 136046 529218 136102
rect 529274 136046 529342 136102
rect 529398 136046 546970 136102
rect 547026 136046 547094 136102
rect 547150 136046 547218 136102
rect 547274 136046 547342 136102
rect 547398 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 39878 135978
rect 39934 135922 40002 135978
rect 40058 135922 70598 135978
rect 70654 135922 70722 135978
rect 70778 135922 101318 135978
rect 101374 135922 101442 135978
rect 101498 135922 132038 135978
rect 132094 135922 132162 135978
rect 132218 135922 162758 135978
rect 162814 135922 162882 135978
rect 162938 135922 193478 135978
rect 193534 135922 193602 135978
rect 193658 135922 224198 135978
rect 224254 135922 224322 135978
rect 224378 135922 254918 135978
rect 254974 135922 255042 135978
rect 255098 135922 285638 135978
rect 285694 135922 285762 135978
rect 285818 135922 316358 135978
rect 316414 135922 316482 135978
rect 316538 135922 347078 135978
rect 347134 135922 347202 135978
rect 347258 135922 377798 135978
rect 377854 135922 377922 135978
rect 377978 135922 408518 135978
rect 408574 135922 408642 135978
rect 408698 135922 439238 135978
rect 439294 135922 439362 135978
rect 439418 135922 469958 135978
rect 470014 135922 470082 135978
rect 470138 135922 500678 135978
rect 500734 135922 500802 135978
rect 500858 135922 528970 135978
rect 529026 135922 529094 135978
rect 529150 135922 529218 135978
rect 529274 135922 529342 135978
rect 529398 135922 546970 135978
rect 547026 135922 547094 135978
rect 547150 135922 547218 135978
rect 547274 135922 547342 135978
rect 547398 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 24518 130350
rect 24574 130294 24642 130350
rect 24698 130294 55238 130350
rect 55294 130294 55362 130350
rect 55418 130294 85958 130350
rect 86014 130294 86082 130350
rect 86138 130294 116678 130350
rect 116734 130294 116802 130350
rect 116858 130294 147398 130350
rect 147454 130294 147522 130350
rect 147578 130294 178118 130350
rect 178174 130294 178242 130350
rect 178298 130294 208838 130350
rect 208894 130294 208962 130350
rect 209018 130294 239558 130350
rect 239614 130294 239682 130350
rect 239738 130294 270278 130350
rect 270334 130294 270402 130350
rect 270458 130294 300998 130350
rect 301054 130294 301122 130350
rect 301178 130294 331718 130350
rect 331774 130294 331842 130350
rect 331898 130294 362438 130350
rect 362494 130294 362562 130350
rect 362618 130294 393158 130350
rect 393214 130294 393282 130350
rect 393338 130294 423878 130350
rect 423934 130294 424002 130350
rect 424058 130294 454598 130350
rect 454654 130294 454722 130350
rect 454778 130294 485318 130350
rect 485374 130294 485442 130350
rect 485498 130294 516038 130350
rect 516094 130294 516162 130350
rect 516218 130294 525250 130350
rect 525306 130294 525374 130350
rect 525430 130294 525498 130350
rect 525554 130294 525622 130350
rect 525678 130294 543250 130350
rect 543306 130294 543374 130350
rect 543430 130294 543498 130350
rect 543554 130294 543622 130350
rect 543678 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 24518 130226
rect 24574 130170 24642 130226
rect 24698 130170 55238 130226
rect 55294 130170 55362 130226
rect 55418 130170 85958 130226
rect 86014 130170 86082 130226
rect 86138 130170 116678 130226
rect 116734 130170 116802 130226
rect 116858 130170 147398 130226
rect 147454 130170 147522 130226
rect 147578 130170 178118 130226
rect 178174 130170 178242 130226
rect 178298 130170 208838 130226
rect 208894 130170 208962 130226
rect 209018 130170 239558 130226
rect 239614 130170 239682 130226
rect 239738 130170 270278 130226
rect 270334 130170 270402 130226
rect 270458 130170 300998 130226
rect 301054 130170 301122 130226
rect 301178 130170 331718 130226
rect 331774 130170 331842 130226
rect 331898 130170 362438 130226
rect 362494 130170 362562 130226
rect 362618 130170 393158 130226
rect 393214 130170 393282 130226
rect 393338 130170 423878 130226
rect 423934 130170 424002 130226
rect 424058 130170 454598 130226
rect 454654 130170 454722 130226
rect 454778 130170 485318 130226
rect 485374 130170 485442 130226
rect 485498 130170 516038 130226
rect 516094 130170 516162 130226
rect 516218 130170 525250 130226
rect 525306 130170 525374 130226
rect 525430 130170 525498 130226
rect 525554 130170 525622 130226
rect 525678 130170 543250 130226
rect 543306 130170 543374 130226
rect 543430 130170 543498 130226
rect 543554 130170 543622 130226
rect 543678 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 24518 130102
rect 24574 130046 24642 130102
rect 24698 130046 55238 130102
rect 55294 130046 55362 130102
rect 55418 130046 85958 130102
rect 86014 130046 86082 130102
rect 86138 130046 116678 130102
rect 116734 130046 116802 130102
rect 116858 130046 147398 130102
rect 147454 130046 147522 130102
rect 147578 130046 178118 130102
rect 178174 130046 178242 130102
rect 178298 130046 208838 130102
rect 208894 130046 208962 130102
rect 209018 130046 239558 130102
rect 239614 130046 239682 130102
rect 239738 130046 270278 130102
rect 270334 130046 270402 130102
rect 270458 130046 300998 130102
rect 301054 130046 301122 130102
rect 301178 130046 331718 130102
rect 331774 130046 331842 130102
rect 331898 130046 362438 130102
rect 362494 130046 362562 130102
rect 362618 130046 393158 130102
rect 393214 130046 393282 130102
rect 393338 130046 423878 130102
rect 423934 130046 424002 130102
rect 424058 130046 454598 130102
rect 454654 130046 454722 130102
rect 454778 130046 485318 130102
rect 485374 130046 485442 130102
rect 485498 130046 516038 130102
rect 516094 130046 516162 130102
rect 516218 130046 525250 130102
rect 525306 130046 525374 130102
rect 525430 130046 525498 130102
rect 525554 130046 525622 130102
rect 525678 130046 543250 130102
rect 543306 130046 543374 130102
rect 543430 130046 543498 130102
rect 543554 130046 543622 130102
rect 543678 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 24518 129978
rect 24574 129922 24642 129978
rect 24698 129922 55238 129978
rect 55294 129922 55362 129978
rect 55418 129922 85958 129978
rect 86014 129922 86082 129978
rect 86138 129922 116678 129978
rect 116734 129922 116802 129978
rect 116858 129922 147398 129978
rect 147454 129922 147522 129978
rect 147578 129922 178118 129978
rect 178174 129922 178242 129978
rect 178298 129922 208838 129978
rect 208894 129922 208962 129978
rect 209018 129922 239558 129978
rect 239614 129922 239682 129978
rect 239738 129922 270278 129978
rect 270334 129922 270402 129978
rect 270458 129922 300998 129978
rect 301054 129922 301122 129978
rect 301178 129922 331718 129978
rect 331774 129922 331842 129978
rect 331898 129922 362438 129978
rect 362494 129922 362562 129978
rect 362618 129922 393158 129978
rect 393214 129922 393282 129978
rect 393338 129922 423878 129978
rect 423934 129922 424002 129978
rect 424058 129922 454598 129978
rect 454654 129922 454722 129978
rect 454778 129922 485318 129978
rect 485374 129922 485442 129978
rect 485498 129922 516038 129978
rect 516094 129922 516162 129978
rect 516218 129922 525250 129978
rect 525306 129922 525374 129978
rect 525430 129922 525498 129978
rect 525554 129922 525622 129978
rect 525678 129922 543250 129978
rect 543306 129922 543374 129978
rect 543430 129922 543498 129978
rect 543554 129922 543622 129978
rect 543678 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 39878 118350
rect 39934 118294 40002 118350
rect 40058 118294 70598 118350
rect 70654 118294 70722 118350
rect 70778 118294 101318 118350
rect 101374 118294 101442 118350
rect 101498 118294 132038 118350
rect 132094 118294 132162 118350
rect 132218 118294 162758 118350
rect 162814 118294 162882 118350
rect 162938 118294 193478 118350
rect 193534 118294 193602 118350
rect 193658 118294 224198 118350
rect 224254 118294 224322 118350
rect 224378 118294 254918 118350
rect 254974 118294 255042 118350
rect 255098 118294 285638 118350
rect 285694 118294 285762 118350
rect 285818 118294 316358 118350
rect 316414 118294 316482 118350
rect 316538 118294 347078 118350
rect 347134 118294 347202 118350
rect 347258 118294 377798 118350
rect 377854 118294 377922 118350
rect 377978 118294 408518 118350
rect 408574 118294 408642 118350
rect 408698 118294 439238 118350
rect 439294 118294 439362 118350
rect 439418 118294 469958 118350
rect 470014 118294 470082 118350
rect 470138 118294 500678 118350
rect 500734 118294 500802 118350
rect 500858 118294 528970 118350
rect 529026 118294 529094 118350
rect 529150 118294 529218 118350
rect 529274 118294 529342 118350
rect 529398 118294 546970 118350
rect 547026 118294 547094 118350
rect 547150 118294 547218 118350
rect 547274 118294 547342 118350
rect 547398 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 39878 118226
rect 39934 118170 40002 118226
rect 40058 118170 70598 118226
rect 70654 118170 70722 118226
rect 70778 118170 101318 118226
rect 101374 118170 101442 118226
rect 101498 118170 132038 118226
rect 132094 118170 132162 118226
rect 132218 118170 162758 118226
rect 162814 118170 162882 118226
rect 162938 118170 193478 118226
rect 193534 118170 193602 118226
rect 193658 118170 224198 118226
rect 224254 118170 224322 118226
rect 224378 118170 254918 118226
rect 254974 118170 255042 118226
rect 255098 118170 285638 118226
rect 285694 118170 285762 118226
rect 285818 118170 316358 118226
rect 316414 118170 316482 118226
rect 316538 118170 347078 118226
rect 347134 118170 347202 118226
rect 347258 118170 377798 118226
rect 377854 118170 377922 118226
rect 377978 118170 408518 118226
rect 408574 118170 408642 118226
rect 408698 118170 439238 118226
rect 439294 118170 439362 118226
rect 439418 118170 469958 118226
rect 470014 118170 470082 118226
rect 470138 118170 500678 118226
rect 500734 118170 500802 118226
rect 500858 118170 528970 118226
rect 529026 118170 529094 118226
rect 529150 118170 529218 118226
rect 529274 118170 529342 118226
rect 529398 118170 546970 118226
rect 547026 118170 547094 118226
rect 547150 118170 547218 118226
rect 547274 118170 547342 118226
rect 547398 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 39878 118102
rect 39934 118046 40002 118102
rect 40058 118046 70598 118102
rect 70654 118046 70722 118102
rect 70778 118046 101318 118102
rect 101374 118046 101442 118102
rect 101498 118046 132038 118102
rect 132094 118046 132162 118102
rect 132218 118046 162758 118102
rect 162814 118046 162882 118102
rect 162938 118046 193478 118102
rect 193534 118046 193602 118102
rect 193658 118046 224198 118102
rect 224254 118046 224322 118102
rect 224378 118046 254918 118102
rect 254974 118046 255042 118102
rect 255098 118046 285638 118102
rect 285694 118046 285762 118102
rect 285818 118046 316358 118102
rect 316414 118046 316482 118102
rect 316538 118046 347078 118102
rect 347134 118046 347202 118102
rect 347258 118046 377798 118102
rect 377854 118046 377922 118102
rect 377978 118046 408518 118102
rect 408574 118046 408642 118102
rect 408698 118046 439238 118102
rect 439294 118046 439362 118102
rect 439418 118046 469958 118102
rect 470014 118046 470082 118102
rect 470138 118046 500678 118102
rect 500734 118046 500802 118102
rect 500858 118046 528970 118102
rect 529026 118046 529094 118102
rect 529150 118046 529218 118102
rect 529274 118046 529342 118102
rect 529398 118046 546970 118102
rect 547026 118046 547094 118102
rect 547150 118046 547218 118102
rect 547274 118046 547342 118102
rect 547398 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 39878 117978
rect 39934 117922 40002 117978
rect 40058 117922 70598 117978
rect 70654 117922 70722 117978
rect 70778 117922 101318 117978
rect 101374 117922 101442 117978
rect 101498 117922 132038 117978
rect 132094 117922 132162 117978
rect 132218 117922 162758 117978
rect 162814 117922 162882 117978
rect 162938 117922 193478 117978
rect 193534 117922 193602 117978
rect 193658 117922 224198 117978
rect 224254 117922 224322 117978
rect 224378 117922 254918 117978
rect 254974 117922 255042 117978
rect 255098 117922 285638 117978
rect 285694 117922 285762 117978
rect 285818 117922 316358 117978
rect 316414 117922 316482 117978
rect 316538 117922 347078 117978
rect 347134 117922 347202 117978
rect 347258 117922 377798 117978
rect 377854 117922 377922 117978
rect 377978 117922 408518 117978
rect 408574 117922 408642 117978
rect 408698 117922 439238 117978
rect 439294 117922 439362 117978
rect 439418 117922 469958 117978
rect 470014 117922 470082 117978
rect 470138 117922 500678 117978
rect 500734 117922 500802 117978
rect 500858 117922 528970 117978
rect 529026 117922 529094 117978
rect 529150 117922 529218 117978
rect 529274 117922 529342 117978
rect 529398 117922 546970 117978
rect 547026 117922 547094 117978
rect 547150 117922 547218 117978
rect 547274 117922 547342 117978
rect 547398 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 24518 112350
rect 24574 112294 24642 112350
rect 24698 112294 55238 112350
rect 55294 112294 55362 112350
rect 55418 112294 85958 112350
rect 86014 112294 86082 112350
rect 86138 112294 116678 112350
rect 116734 112294 116802 112350
rect 116858 112294 147398 112350
rect 147454 112294 147522 112350
rect 147578 112294 178118 112350
rect 178174 112294 178242 112350
rect 178298 112294 208838 112350
rect 208894 112294 208962 112350
rect 209018 112294 239558 112350
rect 239614 112294 239682 112350
rect 239738 112294 270278 112350
rect 270334 112294 270402 112350
rect 270458 112294 300998 112350
rect 301054 112294 301122 112350
rect 301178 112294 331718 112350
rect 331774 112294 331842 112350
rect 331898 112294 362438 112350
rect 362494 112294 362562 112350
rect 362618 112294 393158 112350
rect 393214 112294 393282 112350
rect 393338 112294 423878 112350
rect 423934 112294 424002 112350
rect 424058 112294 454598 112350
rect 454654 112294 454722 112350
rect 454778 112294 485318 112350
rect 485374 112294 485442 112350
rect 485498 112294 516038 112350
rect 516094 112294 516162 112350
rect 516218 112294 525250 112350
rect 525306 112294 525374 112350
rect 525430 112294 525498 112350
rect 525554 112294 525622 112350
rect 525678 112294 543250 112350
rect 543306 112294 543374 112350
rect 543430 112294 543498 112350
rect 543554 112294 543622 112350
rect 543678 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 24518 112226
rect 24574 112170 24642 112226
rect 24698 112170 55238 112226
rect 55294 112170 55362 112226
rect 55418 112170 85958 112226
rect 86014 112170 86082 112226
rect 86138 112170 116678 112226
rect 116734 112170 116802 112226
rect 116858 112170 147398 112226
rect 147454 112170 147522 112226
rect 147578 112170 178118 112226
rect 178174 112170 178242 112226
rect 178298 112170 208838 112226
rect 208894 112170 208962 112226
rect 209018 112170 239558 112226
rect 239614 112170 239682 112226
rect 239738 112170 270278 112226
rect 270334 112170 270402 112226
rect 270458 112170 300998 112226
rect 301054 112170 301122 112226
rect 301178 112170 331718 112226
rect 331774 112170 331842 112226
rect 331898 112170 362438 112226
rect 362494 112170 362562 112226
rect 362618 112170 393158 112226
rect 393214 112170 393282 112226
rect 393338 112170 423878 112226
rect 423934 112170 424002 112226
rect 424058 112170 454598 112226
rect 454654 112170 454722 112226
rect 454778 112170 485318 112226
rect 485374 112170 485442 112226
rect 485498 112170 516038 112226
rect 516094 112170 516162 112226
rect 516218 112170 525250 112226
rect 525306 112170 525374 112226
rect 525430 112170 525498 112226
rect 525554 112170 525622 112226
rect 525678 112170 543250 112226
rect 543306 112170 543374 112226
rect 543430 112170 543498 112226
rect 543554 112170 543622 112226
rect 543678 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 24518 112102
rect 24574 112046 24642 112102
rect 24698 112046 55238 112102
rect 55294 112046 55362 112102
rect 55418 112046 85958 112102
rect 86014 112046 86082 112102
rect 86138 112046 116678 112102
rect 116734 112046 116802 112102
rect 116858 112046 147398 112102
rect 147454 112046 147522 112102
rect 147578 112046 178118 112102
rect 178174 112046 178242 112102
rect 178298 112046 208838 112102
rect 208894 112046 208962 112102
rect 209018 112046 239558 112102
rect 239614 112046 239682 112102
rect 239738 112046 270278 112102
rect 270334 112046 270402 112102
rect 270458 112046 300998 112102
rect 301054 112046 301122 112102
rect 301178 112046 331718 112102
rect 331774 112046 331842 112102
rect 331898 112046 362438 112102
rect 362494 112046 362562 112102
rect 362618 112046 393158 112102
rect 393214 112046 393282 112102
rect 393338 112046 423878 112102
rect 423934 112046 424002 112102
rect 424058 112046 454598 112102
rect 454654 112046 454722 112102
rect 454778 112046 485318 112102
rect 485374 112046 485442 112102
rect 485498 112046 516038 112102
rect 516094 112046 516162 112102
rect 516218 112046 525250 112102
rect 525306 112046 525374 112102
rect 525430 112046 525498 112102
rect 525554 112046 525622 112102
rect 525678 112046 543250 112102
rect 543306 112046 543374 112102
rect 543430 112046 543498 112102
rect 543554 112046 543622 112102
rect 543678 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 24518 111978
rect 24574 111922 24642 111978
rect 24698 111922 55238 111978
rect 55294 111922 55362 111978
rect 55418 111922 85958 111978
rect 86014 111922 86082 111978
rect 86138 111922 116678 111978
rect 116734 111922 116802 111978
rect 116858 111922 147398 111978
rect 147454 111922 147522 111978
rect 147578 111922 178118 111978
rect 178174 111922 178242 111978
rect 178298 111922 208838 111978
rect 208894 111922 208962 111978
rect 209018 111922 239558 111978
rect 239614 111922 239682 111978
rect 239738 111922 270278 111978
rect 270334 111922 270402 111978
rect 270458 111922 300998 111978
rect 301054 111922 301122 111978
rect 301178 111922 331718 111978
rect 331774 111922 331842 111978
rect 331898 111922 362438 111978
rect 362494 111922 362562 111978
rect 362618 111922 393158 111978
rect 393214 111922 393282 111978
rect 393338 111922 423878 111978
rect 423934 111922 424002 111978
rect 424058 111922 454598 111978
rect 454654 111922 454722 111978
rect 454778 111922 485318 111978
rect 485374 111922 485442 111978
rect 485498 111922 516038 111978
rect 516094 111922 516162 111978
rect 516218 111922 525250 111978
rect 525306 111922 525374 111978
rect 525430 111922 525498 111978
rect 525554 111922 525622 111978
rect 525678 111922 543250 111978
rect 543306 111922 543374 111978
rect 543430 111922 543498 111978
rect 543554 111922 543622 111978
rect 543678 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 39878 100350
rect 39934 100294 40002 100350
rect 40058 100294 70598 100350
rect 70654 100294 70722 100350
rect 70778 100294 101318 100350
rect 101374 100294 101442 100350
rect 101498 100294 132038 100350
rect 132094 100294 132162 100350
rect 132218 100294 162758 100350
rect 162814 100294 162882 100350
rect 162938 100294 193478 100350
rect 193534 100294 193602 100350
rect 193658 100294 224198 100350
rect 224254 100294 224322 100350
rect 224378 100294 254918 100350
rect 254974 100294 255042 100350
rect 255098 100294 285638 100350
rect 285694 100294 285762 100350
rect 285818 100294 316358 100350
rect 316414 100294 316482 100350
rect 316538 100294 347078 100350
rect 347134 100294 347202 100350
rect 347258 100294 377798 100350
rect 377854 100294 377922 100350
rect 377978 100294 408518 100350
rect 408574 100294 408642 100350
rect 408698 100294 439238 100350
rect 439294 100294 439362 100350
rect 439418 100294 469958 100350
rect 470014 100294 470082 100350
rect 470138 100294 500678 100350
rect 500734 100294 500802 100350
rect 500858 100294 528970 100350
rect 529026 100294 529094 100350
rect 529150 100294 529218 100350
rect 529274 100294 529342 100350
rect 529398 100294 546970 100350
rect 547026 100294 547094 100350
rect 547150 100294 547218 100350
rect 547274 100294 547342 100350
rect 547398 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 39878 100226
rect 39934 100170 40002 100226
rect 40058 100170 70598 100226
rect 70654 100170 70722 100226
rect 70778 100170 101318 100226
rect 101374 100170 101442 100226
rect 101498 100170 132038 100226
rect 132094 100170 132162 100226
rect 132218 100170 162758 100226
rect 162814 100170 162882 100226
rect 162938 100170 193478 100226
rect 193534 100170 193602 100226
rect 193658 100170 224198 100226
rect 224254 100170 224322 100226
rect 224378 100170 254918 100226
rect 254974 100170 255042 100226
rect 255098 100170 285638 100226
rect 285694 100170 285762 100226
rect 285818 100170 316358 100226
rect 316414 100170 316482 100226
rect 316538 100170 347078 100226
rect 347134 100170 347202 100226
rect 347258 100170 377798 100226
rect 377854 100170 377922 100226
rect 377978 100170 408518 100226
rect 408574 100170 408642 100226
rect 408698 100170 439238 100226
rect 439294 100170 439362 100226
rect 439418 100170 469958 100226
rect 470014 100170 470082 100226
rect 470138 100170 500678 100226
rect 500734 100170 500802 100226
rect 500858 100170 528970 100226
rect 529026 100170 529094 100226
rect 529150 100170 529218 100226
rect 529274 100170 529342 100226
rect 529398 100170 546970 100226
rect 547026 100170 547094 100226
rect 547150 100170 547218 100226
rect 547274 100170 547342 100226
rect 547398 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 39878 100102
rect 39934 100046 40002 100102
rect 40058 100046 70598 100102
rect 70654 100046 70722 100102
rect 70778 100046 101318 100102
rect 101374 100046 101442 100102
rect 101498 100046 132038 100102
rect 132094 100046 132162 100102
rect 132218 100046 162758 100102
rect 162814 100046 162882 100102
rect 162938 100046 193478 100102
rect 193534 100046 193602 100102
rect 193658 100046 224198 100102
rect 224254 100046 224322 100102
rect 224378 100046 254918 100102
rect 254974 100046 255042 100102
rect 255098 100046 285638 100102
rect 285694 100046 285762 100102
rect 285818 100046 316358 100102
rect 316414 100046 316482 100102
rect 316538 100046 347078 100102
rect 347134 100046 347202 100102
rect 347258 100046 377798 100102
rect 377854 100046 377922 100102
rect 377978 100046 408518 100102
rect 408574 100046 408642 100102
rect 408698 100046 439238 100102
rect 439294 100046 439362 100102
rect 439418 100046 469958 100102
rect 470014 100046 470082 100102
rect 470138 100046 500678 100102
rect 500734 100046 500802 100102
rect 500858 100046 528970 100102
rect 529026 100046 529094 100102
rect 529150 100046 529218 100102
rect 529274 100046 529342 100102
rect 529398 100046 546970 100102
rect 547026 100046 547094 100102
rect 547150 100046 547218 100102
rect 547274 100046 547342 100102
rect 547398 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 39878 99978
rect 39934 99922 40002 99978
rect 40058 99922 70598 99978
rect 70654 99922 70722 99978
rect 70778 99922 101318 99978
rect 101374 99922 101442 99978
rect 101498 99922 132038 99978
rect 132094 99922 132162 99978
rect 132218 99922 162758 99978
rect 162814 99922 162882 99978
rect 162938 99922 193478 99978
rect 193534 99922 193602 99978
rect 193658 99922 224198 99978
rect 224254 99922 224322 99978
rect 224378 99922 254918 99978
rect 254974 99922 255042 99978
rect 255098 99922 285638 99978
rect 285694 99922 285762 99978
rect 285818 99922 316358 99978
rect 316414 99922 316482 99978
rect 316538 99922 347078 99978
rect 347134 99922 347202 99978
rect 347258 99922 377798 99978
rect 377854 99922 377922 99978
rect 377978 99922 408518 99978
rect 408574 99922 408642 99978
rect 408698 99922 439238 99978
rect 439294 99922 439362 99978
rect 439418 99922 469958 99978
rect 470014 99922 470082 99978
rect 470138 99922 500678 99978
rect 500734 99922 500802 99978
rect 500858 99922 528970 99978
rect 529026 99922 529094 99978
rect 529150 99922 529218 99978
rect 529274 99922 529342 99978
rect 529398 99922 546970 99978
rect 547026 99922 547094 99978
rect 547150 99922 547218 99978
rect 547274 99922 547342 99978
rect 547398 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 24518 94350
rect 24574 94294 24642 94350
rect 24698 94294 55238 94350
rect 55294 94294 55362 94350
rect 55418 94294 85958 94350
rect 86014 94294 86082 94350
rect 86138 94294 116678 94350
rect 116734 94294 116802 94350
rect 116858 94294 147398 94350
rect 147454 94294 147522 94350
rect 147578 94294 178118 94350
rect 178174 94294 178242 94350
rect 178298 94294 208838 94350
rect 208894 94294 208962 94350
rect 209018 94294 239558 94350
rect 239614 94294 239682 94350
rect 239738 94294 270278 94350
rect 270334 94294 270402 94350
rect 270458 94294 300998 94350
rect 301054 94294 301122 94350
rect 301178 94294 331718 94350
rect 331774 94294 331842 94350
rect 331898 94294 362438 94350
rect 362494 94294 362562 94350
rect 362618 94294 393158 94350
rect 393214 94294 393282 94350
rect 393338 94294 423878 94350
rect 423934 94294 424002 94350
rect 424058 94294 454598 94350
rect 454654 94294 454722 94350
rect 454778 94294 485318 94350
rect 485374 94294 485442 94350
rect 485498 94294 516038 94350
rect 516094 94294 516162 94350
rect 516218 94294 525250 94350
rect 525306 94294 525374 94350
rect 525430 94294 525498 94350
rect 525554 94294 525622 94350
rect 525678 94294 543250 94350
rect 543306 94294 543374 94350
rect 543430 94294 543498 94350
rect 543554 94294 543622 94350
rect 543678 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 24518 94226
rect 24574 94170 24642 94226
rect 24698 94170 55238 94226
rect 55294 94170 55362 94226
rect 55418 94170 85958 94226
rect 86014 94170 86082 94226
rect 86138 94170 116678 94226
rect 116734 94170 116802 94226
rect 116858 94170 147398 94226
rect 147454 94170 147522 94226
rect 147578 94170 178118 94226
rect 178174 94170 178242 94226
rect 178298 94170 208838 94226
rect 208894 94170 208962 94226
rect 209018 94170 239558 94226
rect 239614 94170 239682 94226
rect 239738 94170 270278 94226
rect 270334 94170 270402 94226
rect 270458 94170 300998 94226
rect 301054 94170 301122 94226
rect 301178 94170 331718 94226
rect 331774 94170 331842 94226
rect 331898 94170 362438 94226
rect 362494 94170 362562 94226
rect 362618 94170 393158 94226
rect 393214 94170 393282 94226
rect 393338 94170 423878 94226
rect 423934 94170 424002 94226
rect 424058 94170 454598 94226
rect 454654 94170 454722 94226
rect 454778 94170 485318 94226
rect 485374 94170 485442 94226
rect 485498 94170 516038 94226
rect 516094 94170 516162 94226
rect 516218 94170 525250 94226
rect 525306 94170 525374 94226
rect 525430 94170 525498 94226
rect 525554 94170 525622 94226
rect 525678 94170 543250 94226
rect 543306 94170 543374 94226
rect 543430 94170 543498 94226
rect 543554 94170 543622 94226
rect 543678 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 24518 94102
rect 24574 94046 24642 94102
rect 24698 94046 55238 94102
rect 55294 94046 55362 94102
rect 55418 94046 85958 94102
rect 86014 94046 86082 94102
rect 86138 94046 116678 94102
rect 116734 94046 116802 94102
rect 116858 94046 147398 94102
rect 147454 94046 147522 94102
rect 147578 94046 178118 94102
rect 178174 94046 178242 94102
rect 178298 94046 208838 94102
rect 208894 94046 208962 94102
rect 209018 94046 239558 94102
rect 239614 94046 239682 94102
rect 239738 94046 270278 94102
rect 270334 94046 270402 94102
rect 270458 94046 300998 94102
rect 301054 94046 301122 94102
rect 301178 94046 331718 94102
rect 331774 94046 331842 94102
rect 331898 94046 362438 94102
rect 362494 94046 362562 94102
rect 362618 94046 393158 94102
rect 393214 94046 393282 94102
rect 393338 94046 423878 94102
rect 423934 94046 424002 94102
rect 424058 94046 454598 94102
rect 454654 94046 454722 94102
rect 454778 94046 485318 94102
rect 485374 94046 485442 94102
rect 485498 94046 516038 94102
rect 516094 94046 516162 94102
rect 516218 94046 525250 94102
rect 525306 94046 525374 94102
rect 525430 94046 525498 94102
rect 525554 94046 525622 94102
rect 525678 94046 543250 94102
rect 543306 94046 543374 94102
rect 543430 94046 543498 94102
rect 543554 94046 543622 94102
rect 543678 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 24518 93978
rect 24574 93922 24642 93978
rect 24698 93922 55238 93978
rect 55294 93922 55362 93978
rect 55418 93922 85958 93978
rect 86014 93922 86082 93978
rect 86138 93922 116678 93978
rect 116734 93922 116802 93978
rect 116858 93922 147398 93978
rect 147454 93922 147522 93978
rect 147578 93922 178118 93978
rect 178174 93922 178242 93978
rect 178298 93922 208838 93978
rect 208894 93922 208962 93978
rect 209018 93922 239558 93978
rect 239614 93922 239682 93978
rect 239738 93922 270278 93978
rect 270334 93922 270402 93978
rect 270458 93922 300998 93978
rect 301054 93922 301122 93978
rect 301178 93922 331718 93978
rect 331774 93922 331842 93978
rect 331898 93922 362438 93978
rect 362494 93922 362562 93978
rect 362618 93922 393158 93978
rect 393214 93922 393282 93978
rect 393338 93922 423878 93978
rect 423934 93922 424002 93978
rect 424058 93922 454598 93978
rect 454654 93922 454722 93978
rect 454778 93922 485318 93978
rect 485374 93922 485442 93978
rect 485498 93922 516038 93978
rect 516094 93922 516162 93978
rect 516218 93922 525250 93978
rect 525306 93922 525374 93978
rect 525430 93922 525498 93978
rect 525554 93922 525622 93978
rect 525678 93922 543250 93978
rect 543306 93922 543374 93978
rect 543430 93922 543498 93978
rect 543554 93922 543622 93978
rect 543678 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 39878 82350
rect 39934 82294 40002 82350
rect 40058 82294 70598 82350
rect 70654 82294 70722 82350
rect 70778 82294 101318 82350
rect 101374 82294 101442 82350
rect 101498 82294 132038 82350
rect 132094 82294 132162 82350
rect 132218 82294 162758 82350
rect 162814 82294 162882 82350
rect 162938 82294 193478 82350
rect 193534 82294 193602 82350
rect 193658 82294 224198 82350
rect 224254 82294 224322 82350
rect 224378 82294 254918 82350
rect 254974 82294 255042 82350
rect 255098 82294 285638 82350
rect 285694 82294 285762 82350
rect 285818 82294 316358 82350
rect 316414 82294 316482 82350
rect 316538 82294 347078 82350
rect 347134 82294 347202 82350
rect 347258 82294 377798 82350
rect 377854 82294 377922 82350
rect 377978 82294 408518 82350
rect 408574 82294 408642 82350
rect 408698 82294 439238 82350
rect 439294 82294 439362 82350
rect 439418 82294 469958 82350
rect 470014 82294 470082 82350
rect 470138 82294 500678 82350
rect 500734 82294 500802 82350
rect 500858 82294 528970 82350
rect 529026 82294 529094 82350
rect 529150 82294 529218 82350
rect 529274 82294 529342 82350
rect 529398 82294 546970 82350
rect 547026 82294 547094 82350
rect 547150 82294 547218 82350
rect 547274 82294 547342 82350
rect 547398 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 39878 82226
rect 39934 82170 40002 82226
rect 40058 82170 70598 82226
rect 70654 82170 70722 82226
rect 70778 82170 101318 82226
rect 101374 82170 101442 82226
rect 101498 82170 132038 82226
rect 132094 82170 132162 82226
rect 132218 82170 162758 82226
rect 162814 82170 162882 82226
rect 162938 82170 193478 82226
rect 193534 82170 193602 82226
rect 193658 82170 224198 82226
rect 224254 82170 224322 82226
rect 224378 82170 254918 82226
rect 254974 82170 255042 82226
rect 255098 82170 285638 82226
rect 285694 82170 285762 82226
rect 285818 82170 316358 82226
rect 316414 82170 316482 82226
rect 316538 82170 347078 82226
rect 347134 82170 347202 82226
rect 347258 82170 377798 82226
rect 377854 82170 377922 82226
rect 377978 82170 408518 82226
rect 408574 82170 408642 82226
rect 408698 82170 439238 82226
rect 439294 82170 439362 82226
rect 439418 82170 469958 82226
rect 470014 82170 470082 82226
rect 470138 82170 500678 82226
rect 500734 82170 500802 82226
rect 500858 82170 528970 82226
rect 529026 82170 529094 82226
rect 529150 82170 529218 82226
rect 529274 82170 529342 82226
rect 529398 82170 546970 82226
rect 547026 82170 547094 82226
rect 547150 82170 547218 82226
rect 547274 82170 547342 82226
rect 547398 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 39878 82102
rect 39934 82046 40002 82102
rect 40058 82046 70598 82102
rect 70654 82046 70722 82102
rect 70778 82046 101318 82102
rect 101374 82046 101442 82102
rect 101498 82046 132038 82102
rect 132094 82046 132162 82102
rect 132218 82046 162758 82102
rect 162814 82046 162882 82102
rect 162938 82046 193478 82102
rect 193534 82046 193602 82102
rect 193658 82046 224198 82102
rect 224254 82046 224322 82102
rect 224378 82046 254918 82102
rect 254974 82046 255042 82102
rect 255098 82046 285638 82102
rect 285694 82046 285762 82102
rect 285818 82046 316358 82102
rect 316414 82046 316482 82102
rect 316538 82046 347078 82102
rect 347134 82046 347202 82102
rect 347258 82046 377798 82102
rect 377854 82046 377922 82102
rect 377978 82046 408518 82102
rect 408574 82046 408642 82102
rect 408698 82046 439238 82102
rect 439294 82046 439362 82102
rect 439418 82046 469958 82102
rect 470014 82046 470082 82102
rect 470138 82046 500678 82102
rect 500734 82046 500802 82102
rect 500858 82046 528970 82102
rect 529026 82046 529094 82102
rect 529150 82046 529218 82102
rect 529274 82046 529342 82102
rect 529398 82046 546970 82102
rect 547026 82046 547094 82102
rect 547150 82046 547218 82102
rect 547274 82046 547342 82102
rect 547398 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 39878 81978
rect 39934 81922 40002 81978
rect 40058 81922 70598 81978
rect 70654 81922 70722 81978
rect 70778 81922 101318 81978
rect 101374 81922 101442 81978
rect 101498 81922 132038 81978
rect 132094 81922 132162 81978
rect 132218 81922 162758 81978
rect 162814 81922 162882 81978
rect 162938 81922 193478 81978
rect 193534 81922 193602 81978
rect 193658 81922 224198 81978
rect 224254 81922 224322 81978
rect 224378 81922 254918 81978
rect 254974 81922 255042 81978
rect 255098 81922 285638 81978
rect 285694 81922 285762 81978
rect 285818 81922 316358 81978
rect 316414 81922 316482 81978
rect 316538 81922 347078 81978
rect 347134 81922 347202 81978
rect 347258 81922 377798 81978
rect 377854 81922 377922 81978
rect 377978 81922 408518 81978
rect 408574 81922 408642 81978
rect 408698 81922 439238 81978
rect 439294 81922 439362 81978
rect 439418 81922 469958 81978
rect 470014 81922 470082 81978
rect 470138 81922 500678 81978
rect 500734 81922 500802 81978
rect 500858 81922 528970 81978
rect 529026 81922 529094 81978
rect 529150 81922 529218 81978
rect 529274 81922 529342 81978
rect 529398 81922 546970 81978
rect 547026 81922 547094 81978
rect 547150 81922 547218 81978
rect 547274 81922 547342 81978
rect 547398 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 24518 76350
rect 24574 76294 24642 76350
rect 24698 76294 55238 76350
rect 55294 76294 55362 76350
rect 55418 76294 85958 76350
rect 86014 76294 86082 76350
rect 86138 76294 116678 76350
rect 116734 76294 116802 76350
rect 116858 76294 147398 76350
rect 147454 76294 147522 76350
rect 147578 76294 178118 76350
rect 178174 76294 178242 76350
rect 178298 76294 208838 76350
rect 208894 76294 208962 76350
rect 209018 76294 239558 76350
rect 239614 76294 239682 76350
rect 239738 76294 270278 76350
rect 270334 76294 270402 76350
rect 270458 76294 300998 76350
rect 301054 76294 301122 76350
rect 301178 76294 331718 76350
rect 331774 76294 331842 76350
rect 331898 76294 362438 76350
rect 362494 76294 362562 76350
rect 362618 76294 393158 76350
rect 393214 76294 393282 76350
rect 393338 76294 423878 76350
rect 423934 76294 424002 76350
rect 424058 76294 454598 76350
rect 454654 76294 454722 76350
rect 454778 76294 485318 76350
rect 485374 76294 485442 76350
rect 485498 76294 516038 76350
rect 516094 76294 516162 76350
rect 516218 76294 525250 76350
rect 525306 76294 525374 76350
rect 525430 76294 525498 76350
rect 525554 76294 525622 76350
rect 525678 76294 543250 76350
rect 543306 76294 543374 76350
rect 543430 76294 543498 76350
rect 543554 76294 543622 76350
rect 543678 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 24518 76226
rect 24574 76170 24642 76226
rect 24698 76170 55238 76226
rect 55294 76170 55362 76226
rect 55418 76170 85958 76226
rect 86014 76170 86082 76226
rect 86138 76170 116678 76226
rect 116734 76170 116802 76226
rect 116858 76170 147398 76226
rect 147454 76170 147522 76226
rect 147578 76170 178118 76226
rect 178174 76170 178242 76226
rect 178298 76170 208838 76226
rect 208894 76170 208962 76226
rect 209018 76170 239558 76226
rect 239614 76170 239682 76226
rect 239738 76170 270278 76226
rect 270334 76170 270402 76226
rect 270458 76170 300998 76226
rect 301054 76170 301122 76226
rect 301178 76170 331718 76226
rect 331774 76170 331842 76226
rect 331898 76170 362438 76226
rect 362494 76170 362562 76226
rect 362618 76170 393158 76226
rect 393214 76170 393282 76226
rect 393338 76170 423878 76226
rect 423934 76170 424002 76226
rect 424058 76170 454598 76226
rect 454654 76170 454722 76226
rect 454778 76170 485318 76226
rect 485374 76170 485442 76226
rect 485498 76170 516038 76226
rect 516094 76170 516162 76226
rect 516218 76170 525250 76226
rect 525306 76170 525374 76226
rect 525430 76170 525498 76226
rect 525554 76170 525622 76226
rect 525678 76170 543250 76226
rect 543306 76170 543374 76226
rect 543430 76170 543498 76226
rect 543554 76170 543622 76226
rect 543678 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 24518 76102
rect 24574 76046 24642 76102
rect 24698 76046 55238 76102
rect 55294 76046 55362 76102
rect 55418 76046 85958 76102
rect 86014 76046 86082 76102
rect 86138 76046 116678 76102
rect 116734 76046 116802 76102
rect 116858 76046 147398 76102
rect 147454 76046 147522 76102
rect 147578 76046 178118 76102
rect 178174 76046 178242 76102
rect 178298 76046 208838 76102
rect 208894 76046 208962 76102
rect 209018 76046 239558 76102
rect 239614 76046 239682 76102
rect 239738 76046 270278 76102
rect 270334 76046 270402 76102
rect 270458 76046 300998 76102
rect 301054 76046 301122 76102
rect 301178 76046 331718 76102
rect 331774 76046 331842 76102
rect 331898 76046 362438 76102
rect 362494 76046 362562 76102
rect 362618 76046 393158 76102
rect 393214 76046 393282 76102
rect 393338 76046 423878 76102
rect 423934 76046 424002 76102
rect 424058 76046 454598 76102
rect 454654 76046 454722 76102
rect 454778 76046 485318 76102
rect 485374 76046 485442 76102
rect 485498 76046 516038 76102
rect 516094 76046 516162 76102
rect 516218 76046 525250 76102
rect 525306 76046 525374 76102
rect 525430 76046 525498 76102
rect 525554 76046 525622 76102
rect 525678 76046 543250 76102
rect 543306 76046 543374 76102
rect 543430 76046 543498 76102
rect 543554 76046 543622 76102
rect 543678 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 24518 75978
rect 24574 75922 24642 75978
rect 24698 75922 55238 75978
rect 55294 75922 55362 75978
rect 55418 75922 85958 75978
rect 86014 75922 86082 75978
rect 86138 75922 116678 75978
rect 116734 75922 116802 75978
rect 116858 75922 147398 75978
rect 147454 75922 147522 75978
rect 147578 75922 178118 75978
rect 178174 75922 178242 75978
rect 178298 75922 208838 75978
rect 208894 75922 208962 75978
rect 209018 75922 239558 75978
rect 239614 75922 239682 75978
rect 239738 75922 270278 75978
rect 270334 75922 270402 75978
rect 270458 75922 300998 75978
rect 301054 75922 301122 75978
rect 301178 75922 331718 75978
rect 331774 75922 331842 75978
rect 331898 75922 362438 75978
rect 362494 75922 362562 75978
rect 362618 75922 393158 75978
rect 393214 75922 393282 75978
rect 393338 75922 423878 75978
rect 423934 75922 424002 75978
rect 424058 75922 454598 75978
rect 454654 75922 454722 75978
rect 454778 75922 485318 75978
rect 485374 75922 485442 75978
rect 485498 75922 516038 75978
rect 516094 75922 516162 75978
rect 516218 75922 525250 75978
rect 525306 75922 525374 75978
rect 525430 75922 525498 75978
rect 525554 75922 525622 75978
rect 525678 75922 543250 75978
rect 543306 75922 543374 75978
rect 543430 75922 543498 75978
rect 543554 75922 543622 75978
rect 543678 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 39878 64350
rect 39934 64294 40002 64350
rect 40058 64294 70598 64350
rect 70654 64294 70722 64350
rect 70778 64294 101318 64350
rect 101374 64294 101442 64350
rect 101498 64294 132038 64350
rect 132094 64294 132162 64350
rect 132218 64294 162758 64350
rect 162814 64294 162882 64350
rect 162938 64294 193478 64350
rect 193534 64294 193602 64350
rect 193658 64294 224198 64350
rect 224254 64294 224322 64350
rect 224378 64294 254918 64350
rect 254974 64294 255042 64350
rect 255098 64294 285638 64350
rect 285694 64294 285762 64350
rect 285818 64294 316358 64350
rect 316414 64294 316482 64350
rect 316538 64294 347078 64350
rect 347134 64294 347202 64350
rect 347258 64294 377798 64350
rect 377854 64294 377922 64350
rect 377978 64294 408518 64350
rect 408574 64294 408642 64350
rect 408698 64294 439238 64350
rect 439294 64294 439362 64350
rect 439418 64294 469958 64350
rect 470014 64294 470082 64350
rect 470138 64294 500678 64350
rect 500734 64294 500802 64350
rect 500858 64294 528970 64350
rect 529026 64294 529094 64350
rect 529150 64294 529218 64350
rect 529274 64294 529342 64350
rect 529398 64294 546970 64350
rect 547026 64294 547094 64350
rect 547150 64294 547218 64350
rect 547274 64294 547342 64350
rect 547398 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 39878 64226
rect 39934 64170 40002 64226
rect 40058 64170 70598 64226
rect 70654 64170 70722 64226
rect 70778 64170 101318 64226
rect 101374 64170 101442 64226
rect 101498 64170 132038 64226
rect 132094 64170 132162 64226
rect 132218 64170 162758 64226
rect 162814 64170 162882 64226
rect 162938 64170 193478 64226
rect 193534 64170 193602 64226
rect 193658 64170 224198 64226
rect 224254 64170 224322 64226
rect 224378 64170 254918 64226
rect 254974 64170 255042 64226
rect 255098 64170 285638 64226
rect 285694 64170 285762 64226
rect 285818 64170 316358 64226
rect 316414 64170 316482 64226
rect 316538 64170 347078 64226
rect 347134 64170 347202 64226
rect 347258 64170 377798 64226
rect 377854 64170 377922 64226
rect 377978 64170 408518 64226
rect 408574 64170 408642 64226
rect 408698 64170 439238 64226
rect 439294 64170 439362 64226
rect 439418 64170 469958 64226
rect 470014 64170 470082 64226
rect 470138 64170 500678 64226
rect 500734 64170 500802 64226
rect 500858 64170 528970 64226
rect 529026 64170 529094 64226
rect 529150 64170 529218 64226
rect 529274 64170 529342 64226
rect 529398 64170 546970 64226
rect 547026 64170 547094 64226
rect 547150 64170 547218 64226
rect 547274 64170 547342 64226
rect 547398 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 39878 64102
rect 39934 64046 40002 64102
rect 40058 64046 70598 64102
rect 70654 64046 70722 64102
rect 70778 64046 101318 64102
rect 101374 64046 101442 64102
rect 101498 64046 132038 64102
rect 132094 64046 132162 64102
rect 132218 64046 162758 64102
rect 162814 64046 162882 64102
rect 162938 64046 193478 64102
rect 193534 64046 193602 64102
rect 193658 64046 224198 64102
rect 224254 64046 224322 64102
rect 224378 64046 254918 64102
rect 254974 64046 255042 64102
rect 255098 64046 285638 64102
rect 285694 64046 285762 64102
rect 285818 64046 316358 64102
rect 316414 64046 316482 64102
rect 316538 64046 347078 64102
rect 347134 64046 347202 64102
rect 347258 64046 377798 64102
rect 377854 64046 377922 64102
rect 377978 64046 408518 64102
rect 408574 64046 408642 64102
rect 408698 64046 439238 64102
rect 439294 64046 439362 64102
rect 439418 64046 469958 64102
rect 470014 64046 470082 64102
rect 470138 64046 500678 64102
rect 500734 64046 500802 64102
rect 500858 64046 528970 64102
rect 529026 64046 529094 64102
rect 529150 64046 529218 64102
rect 529274 64046 529342 64102
rect 529398 64046 546970 64102
rect 547026 64046 547094 64102
rect 547150 64046 547218 64102
rect 547274 64046 547342 64102
rect 547398 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 39878 63978
rect 39934 63922 40002 63978
rect 40058 63922 70598 63978
rect 70654 63922 70722 63978
rect 70778 63922 101318 63978
rect 101374 63922 101442 63978
rect 101498 63922 132038 63978
rect 132094 63922 132162 63978
rect 132218 63922 162758 63978
rect 162814 63922 162882 63978
rect 162938 63922 193478 63978
rect 193534 63922 193602 63978
rect 193658 63922 224198 63978
rect 224254 63922 224322 63978
rect 224378 63922 254918 63978
rect 254974 63922 255042 63978
rect 255098 63922 285638 63978
rect 285694 63922 285762 63978
rect 285818 63922 316358 63978
rect 316414 63922 316482 63978
rect 316538 63922 347078 63978
rect 347134 63922 347202 63978
rect 347258 63922 377798 63978
rect 377854 63922 377922 63978
rect 377978 63922 408518 63978
rect 408574 63922 408642 63978
rect 408698 63922 439238 63978
rect 439294 63922 439362 63978
rect 439418 63922 469958 63978
rect 470014 63922 470082 63978
rect 470138 63922 500678 63978
rect 500734 63922 500802 63978
rect 500858 63922 528970 63978
rect 529026 63922 529094 63978
rect 529150 63922 529218 63978
rect 529274 63922 529342 63978
rect 529398 63922 546970 63978
rect 547026 63922 547094 63978
rect 547150 63922 547218 63978
rect 547274 63922 547342 63978
rect 547398 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 24518 58350
rect 24574 58294 24642 58350
rect 24698 58294 55238 58350
rect 55294 58294 55362 58350
rect 55418 58294 85958 58350
rect 86014 58294 86082 58350
rect 86138 58294 116678 58350
rect 116734 58294 116802 58350
rect 116858 58294 147398 58350
rect 147454 58294 147522 58350
rect 147578 58294 178118 58350
rect 178174 58294 178242 58350
rect 178298 58294 208838 58350
rect 208894 58294 208962 58350
rect 209018 58294 239558 58350
rect 239614 58294 239682 58350
rect 239738 58294 270278 58350
rect 270334 58294 270402 58350
rect 270458 58294 300998 58350
rect 301054 58294 301122 58350
rect 301178 58294 331718 58350
rect 331774 58294 331842 58350
rect 331898 58294 362438 58350
rect 362494 58294 362562 58350
rect 362618 58294 393158 58350
rect 393214 58294 393282 58350
rect 393338 58294 423878 58350
rect 423934 58294 424002 58350
rect 424058 58294 454598 58350
rect 454654 58294 454722 58350
rect 454778 58294 485318 58350
rect 485374 58294 485442 58350
rect 485498 58294 516038 58350
rect 516094 58294 516162 58350
rect 516218 58294 525250 58350
rect 525306 58294 525374 58350
rect 525430 58294 525498 58350
rect 525554 58294 525622 58350
rect 525678 58294 543250 58350
rect 543306 58294 543374 58350
rect 543430 58294 543498 58350
rect 543554 58294 543622 58350
rect 543678 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 24518 58226
rect 24574 58170 24642 58226
rect 24698 58170 55238 58226
rect 55294 58170 55362 58226
rect 55418 58170 85958 58226
rect 86014 58170 86082 58226
rect 86138 58170 116678 58226
rect 116734 58170 116802 58226
rect 116858 58170 147398 58226
rect 147454 58170 147522 58226
rect 147578 58170 178118 58226
rect 178174 58170 178242 58226
rect 178298 58170 208838 58226
rect 208894 58170 208962 58226
rect 209018 58170 239558 58226
rect 239614 58170 239682 58226
rect 239738 58170 270278 58226
rect 270334 58170 270402 58226
rect 270458 58170 300998 58226
rect 301054 58170 301122 58226
rect 301178 58170 331718 58226
rect 331774 58170 331842 58226
rect 331898 58170 362438 58226
rect 362494 58170 362562 58226
rect 362618 58170 393158 58226
rect 393214 58170 393282 58226
rect 393338 58170 423878 58226
rect 423934 58170 424002 58226
rect 424058 58170 454598 58226
rect 454654 58170 454722 58226
rect 454778 58170 485318 58226
rect 485374 58170 485442 58226
rect 485498 58170 516038 58226
rect 516094 58170 516162 58226
rect 516218 58170 525250 58226
rect 525306 58170 525374 58226
rect 525430 58170 525498 58226
rect 525554 58170 525622 58226
rect 525678 58170 543250 58226
rect 543306 58170 543374 58226
rect 543430 58170 543498 58226
rect 543554 58170 543622 58226
rect 543678 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 24518 58102
rect 24574 58046 24642 58102
rect 24698 58046 55238 58102
rect 55294 58046 55362 58102
rect 55418 58046 85958 58102
rect 86014 58046 86082 58102
rect 86138 58046 116678 58102
rect 116734 58046 116802 58102
rect 116858 58046 147398 58102
rect 147454 58046 147522 58102
rect 147578 58046 178118 58102
rect 178174 58046 178242 58102
rect 178298 58046 208838 58102
rect 208894 58046 208962 58102
rect 209018 58046 239558 58102
rect 239614 58046 239682 58102
rect 239738 58046 270278 58102
rect 270334 58046 270402 58102
rect 270458 58046 300998 58102
rect 301054 58046 301122 58102
rect 301178 58046 331718 58102
rect 331774 58046 331842 58102
rect 331898 58046 362438 58102
rect 362494 58046 362562 58102
rect 362618 58046 393158 58102
rect 393214 58046 393282 58102
rect 393338 58046 423878 58102
rect 423934 58046 424002 58102
rect 424058 58046 454598 58102
rect 454654 58046 454722 58102
rect 454778 58046 485318 58102
rect 485374 58046 485442 58102
rect 485498 58046 516038 58102
rect 516094 58046 516162 58102
rect 516218 58046 525250 58102
rect 525306 58046 525374 58102
rect 525430 58046 525498 58102
rect 525554 58046 525622 58102
rect 525678 58046 543250 58102
rect 543306 58046 543374 58102
rect 543430 58046 543498 58102
rect 543554 58046 543622 58102
rect 543678 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 24518 57978
rect 24574 57922 24642 57978
rect 24698 57922 55238 57978
rect 55294 57922 55362 57978
rect 55418 57922 85958 57978
rect 86014 57922 86082 57978
rect 86138 57922 116678 57978
rect 116734 57922 116802 57978
rect 116858 57922 147398 57978
rect 147454 57922 147522 57978
rect 147578 57922 178118 57978
rect 178174 57922 178242 57978
rect 178298 57922 208838 57978
rect 208894 57922 208962 57978
rect 209018 57922 239558 57978
rect 239614 57922 239682 57978
rect 239738 57922 270278 57978
rect 270334 57922 270402 57978
rect 270458 57922 300998 57978
rect 301054 57922 301122 57978
rect 301178 57922 331718 57978
rect 331774 57922 331842 57978
rect 331898 57922 362438 57978
rect 362494 57922 362562 57978
rect 362618 57922 393158 57978
rect 393214 57922 393282 57978
rect 393338 57922 423878 57978
rect 423934 57922 424002 57978
rect 424058 57922 454598 57978
rect 454654 57922 454722 57978
rect 454778 57922 485318 57978
rect 485374 57922 485442 57978
rect 485498 57922 516038 57978
rect 516094 57922 516162 57978
rect 516218 57922 525250 57978
rect 525306 57922 525374 57978
rect 525430 57922 525498 57978
rect 525554 57922 525622 57978
rect 525678 57922 543250 57978
rect 543306 57922 543374 57978
rect 543430 57922 543498 57978
rect 543554 57922 543622 57978
rect 543678 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 39878 46350
rect 39934 46294 40002 46350
rect 40058 46294 70598 46350
rect 70654 46294 70722 46350
rect 70778 46294 101318 46350
rect 101374 46294 101442 46350
rect 101498 46294 132038 46350
rect 132094 46294 132162 46350
rect 132218 46294 162758 46350
rect 162814 46294 162882 46350
rect 162938 46294 193478 46350
rect 193534 46294 193602 46350
rect 193658 46294 224198 46350
rect 224254 46294 224322 46350
rect 224378 46294 254918 46350
rect 254974 46294 255042 46350
rect 255098 46294 285638 46350
rect 285694 46294 285762 46350
rect 285818 46294 316358 46350
rect 316414 46294 316482 46350
rect 316538 46294 347078 46350
rect 347134 46294 347202 46350
rect 347258 46294 377798 46350
rect 377854 46294 377922 46350
rect 377978 46294 408518 46350
rect 408574 46294 408642 46350
rect 408698 46294 439238 46350
rect 439294 46294 439362 46350
rect 439418 46294 469958 46350
rect 470014 46294 470082 46350
rect 470138 46294 500678 46350
rect 500734 46294 500802 46350
rect 500858 46294 528970 46350
rect 529026 46294 529094 46350
rect 529150 46294 529218 46350
rect 529274 46294 529342 46350
rect 529398 46294 546970 46350
rect 547026 46294 547094 46350
rect 547150 46294 547218 46350
rect 547274 46294 547342 46350
rect 547398 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 39878 46226
rect 39934 46170 40002 46226
rect 40058 46170 70598 46226
rect 70654 46170 70722 46226
rect 70778 46170 101318 46226
rect 101374 46170 101442 46226
rect 101498 46170 132038 46226
rect 132094 46170 132162 46226
rect 132218 46170 162758 46226
rect 162814 46170 162882 46226
rect 162938 46170 193478 46226
rect 193534 46170 193602 46226
rect 193658 46170 224198 46226
rect 224254 46170 224322 46226
rect 224378 46170 254918 46226
rect 254974 46170 255042 46226
rect 255098 46170 285638 46226
rect 285694 46170 285762 46226
rect 285818 46170 316358 46226
rect 316414 46170 316482 46226
rect 316538 46170 347078 46226
rect 347134 46170 347202 46226
rect 347258 46170 377798 46226
rect 377854 46170 377922 46226
rect 377978 46170 408518 46226
rect 408574 46170 408642 46226
rect 408698 46170 439238 46226
rect 439294 46170 439362 46226
rect 439418 46170 469958 46226
rect 470014 46170 470082 46226
rect 470138 46170 500678 46226
rect 500734 46170 500802 46226
rect 500858 46170 528970 46226
rect 529026 46170 529094 46226
rect 529150 46170 529218 46226
rect 529274 46170 529342 46226
rect 529398 46170 546970 46226
rect 547026 46170 547094 46226
rect 547150 46170 547218 46226
rect 547274 46170 547342 46226
rect 547398 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 39878 46102
rect 39934 46046 40002 46102
rect 40058 46046 70598 46102
rect 70654 46046 70722 46102
rect 70778 46046 101318 46102
rect 101374 46046 101442 46102
rect 101498 46046 132038 46102
rect 132094 46046 132162 46102
rect 132218 46046 162758 46102
rect 162814 46046 162882 46102
rect 162938 46046 193478 46102
rect 193534 46046 193602 46102
rect 193658 46046 224198 46102
rect 224254 46046 224322 46102
rect 224378 46046 254918 46102
rect 254974 46046 255042 46102
rect 255098 46046 285638 46102
rect 285694 46046 285762 46102
rect 285818 46046 316358 46102
rect 316414 46046 316482 46102
rect 316538 46046 347078 46102
rect 347134 46046 347202 46102
rect 347258 46046 377798 46102
rect 377854 46046 377922 46102
rect 377978 46046 408518 46102
rect 408574 46046 408642 46102
rect 408698 46046 439238 46102
rect 439294 46046 439362 46102
rect 439418 46046 469958 46102
rect 470014 46046 470082 46102
rect 470138 46046 500678 46102
rect 500734 46046 500802 46102
rect 500858 46046 528970 46102
rect 529026 46046 529094 46102
rect 529150 46046 529218 46102
rect 529274 46046 529342 46102
rect 529398 46046 546970 46102
rect 547026 46046 547094 46102
rect 547150 46046 547218 46102
rect 547274 46046 547342 46102
rect 547398 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 39878 45978
rect 39934 45922 40002 45978
rect 40058 45922 70598 45978
rect 70654 45922 70722 45978
rect 70778 45922 101318 45978
rect 101374 45922 101442 45978
rect 101498 45922 132038 45978
rect 132094 45922 132162 45978
rect 132218 45922 162758 45978
rect 162814 45922 162882 45978
rect 162938 45922 193478 45978
rect 193534 45922 193602 45978
rect 193658 45922 224198 45978
rect 224254 45922 224322 45978
rect 224378 45922 254918 45978
rect 254974 45922 255042 45978
rect 255098 45922 285638 45978
rect 285694 45922 285762 45978
rect 285818 45922 316358 45978
rect 316414 45922 316482 45978
rect 316538 45922 347078 45978
rect 347134 45922 347202 45978
rect 347258 45922 377798 45978
rect 377854 45922 377922 45978
rect 377978 45922 408518 45978
rect 408574 45922 408642 45978
rect 408698 45922 439238 45978
rect 439294 45922 439362 45978
rect 439418 45922 469958 45978
rect 470014 45922 470082 45978
rect 470138 45922 500678 45978
rect 500734 45922 500802 45978
rect 500858 45922 528970 45978
rect 529026 45922 529094 45978
rect 529150 45922 529218 45978
rect 529274 45922 529342 45978
rect 529398 45922 546970 45978
rect 547026 45922 547094 45978
rect 547150 45922 547218 45978
rect 547274 45922 547342 45978
rect 547398 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 24518 40350
rect 24574 40294 24642 40350
rect 24698 40294 55238 40350
rect 55294 40294 55362 40350
rect 55418 40294 85958 40350
rect 86014 40294 86082 40350
rect 86138 40294 116678 40350
rect 116734 40294 116802 40350
rect 116858 40294 147398 40350
rect 147454 40294 147522 40350
rect 147578 40294 178118 40350
rect 178174 40294 178242 40350
rect 178298 40294 208838 40350
rect 208894 40294 208962 40350
rect 209018 40294 239558 40350
rect 239614 40294 239682 40350
rect 239738 40294 270278 40350
rect 270334 40294 270402 40350
rect 270458 40294 300998 40350
rect 301054 40294 301122 40350
rect 301178 40294 331718 40350
rect 331774 40294 331842 40350
rect 331898 40294 362438 40350
rect 362494 40294 362562 40350
rect 362618 40294 393158 40350
rect 393214 40294 393282 40350
rect 393338 40294 423878 40350
rect 423934 40294 424002 40350
rect 424058 40294 454598 40350
rect 454654 40294 454722 40350
rect 454778 40294 485318 40350
rect 485374 40294 485442 40350
rect 485498 40294 516038 40350
rect 516094 40294 516162 40350
rect 516218 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 24518 40226
rect 24574 40170 24642 40226
rect 24698 40170 55238 40226
rect 55294 40170 55362 40226
rect 55418 40170 85958 40226
rect 86014 40170 86082 40226
rect 86138 40170 116678 40226
rect 116734 40170 116802 40226
rect 116858 40170 147398 40226
rect 147454 40170 147522 40226
rect 147578 40170 178118 40226
rect 178174 40170 178242 40226
rect 178298 40170 208838 40226
rect 208894 40170 208962 40226
rect 209018 40170 239558 40226
rect 239614 40170 239682 40226
rect 239738 40170 270278 40226
rect 270334 40170 270402 40226
rect 270458 40170 300998 40226
rect 301054 40170 301122 40226
rect 301178 40170 331718 40226
rect 331774 40170 331842 40226
rect 331898 40170 362438 40226
rect 362494 40170 362562 40226
rect 362618 40170 393158 40226
rect 393214 40170 393282 40226
rect 393338 40170 423878 40226
rect 423934 40170 424002 40226
rect 424058 40170 454598 40226
rect 454654 40170 454722 40226
rect 454778 40170 485318 40226
rect 485374 40170 485442 40226
rect 485498 40170 516038 40226
rect 516094 40170 516162 40226
rect 516218 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 24518 40102
rect 24574 40046 24642 40102
rect 24698 40046 55238 40102
rect 55294 40046 55362 40102
rect 55418 40046 85958 40102
rect 86014 40046 86082 40102
rect 86138 40046 116678 40102
rect 116734 40046 116802 40102
rect 116858 40046 147398 40102
rect 147454 40046 147522 40102
rect 147578 40046 178118 40102
rect 178174 40046 178242 40102
rect 178298 40046 208838 40102
rect 208894 40046 208962 40102
rect 209018 40046 239558 40102
rect 239614 40046 239682 40102
rect 239738 40046 270278 40102
rect 270334 40046 270402 40102
rect 270458 40046 300998 40102
rect 301054 40046 301122 40102
rect 301178 40046 331718 40102
rect 331774 40046 331842 40102
rect 331898 40046 362438 40102
rect 362494 40046 362562 40102
rect 362618 40046 393158 40102
rect 393214 40046 393282 40102
rect 393338 40046 423878 40102
rect 423934 40046 424002 40102
rect 424058 40046 454598 40102
rect 454654 40046 454722 40102
rect 454778 40046 485318 40102
rect 485374 40046 485442 40102
rect 485498 40046 516038 40102
rect 516094 40046 516162 40102
rect 516218 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 24518 39978
rect 24574 39922 24642 39978
rect 24698 39922 55238 39978
rect 55294 39922 55362 39978
rect 55418 39922 85958 39978
rect 86014 39922 86082 39978
rect 86138 39922 116678 39978
rect 116734 39922 116802 39978
rect 116858 39922 147398 39978
rect 147454 39922 147522 39978
rect 147578 39922 178118 39978
rect 178174 39922 178242 39978
rect 178298 39922 208838 39978
rect 208894 39922 208962 39978
rect 209018 39922 239558 39978
rect 239614 39922 239682 39978
rect 239738 39922 270278 39978
rect 270334 39922 270402 39978
rect 270458 39922 300998 39978
rect 301054 39922 301122 39978
rect 301178 39922 331718 39978
rect 331774 39922 331842 39978
rect 331898 39922 362438 39978
rect 362494 39922 362562 39978
rect 362618 39922 393158 39978
rect 393214 39922 393282 39978
rect 393338 39922 423878 39978
rect 423934 39922 424002 39978
rect 424058 39922 454598 39978
rect 454654 39922 454722 39978
rect 454778 39922 485318 39978
rect 485374 39922 485442 39978
rect 485498 39922 516038 39978
rect 516094 39922 516162 39978
rect 516218 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 39878 28350
rect 39934 28294 40002 28350
rect 40058 28294 70598 28350
rect 70654 28294 70722 28350
rect 70778 28294 101318 28350
rect 101374 28294 101442 28350
rect 101498 28294 132038 28350
rect 132094 28294 132162 28350
rect 132218 28294 162758 28350
rect 162814 28294 162882 28350
rect 162938 28294 193478 28350
rect 193534 28294 193602 28350
rect 193658 28294 224198 28350
rect 224254 28294 224322 28350
rect 224378 28294 254918 28350
rect 254974 28294 255042 28350
rect 255098 28294 285638 28350
rect 285694 28294 285762 28350
rect 285818 28294 316358 28350
rect 316414 28294 316482 28350
rect 316538 28294 347078 28350
rect 347134 28294 347202 28350
rect 347258 28294 377798 28350
rect 377854 28294 377922 28350
rect 377978 28294 408518 28350
rect 408574 28294 408642 28350
rect 408698 28294 439238 28350
rect 439294 28294 439362 28350
rect 439418 28294 469958 28350
rect 470014 28294 470082 28350
rect 470138 28294 500678 28350
rect 500734 28294 500802 28350
rect 500858 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 39878 28226
rect 39934 28170 40002 28226
rect 40058 28170 70598 28226
rect 70654 28170 70722 28226
rect 70778 28170 101318 28226
rect 101374 28170 101442 28226
rect 101498 28170 132038 28226
rect 132094 28170 132162 28226
rect 132218 28170 162758 28226
rect 162814 28170 162882 28226
rect 162938 28170 193478 28226
rect 193534 28170 193602 28226
rect 193658 28170 224198 28226
rect 224254 28170 224322 28226
rect 224378 28170 254918 28226
rect 254974 28170 255042 28226
rect 255098 28170 285638 28226
rect 285694 28170 285762 28226
rect 285818 28170 316358 28226
rect 316414 28170 316482 28226
rect 316538 28170 347078 28226
rect 347134 28170 347202 28226
rect 347258 28170 377798 28226
rect 377854 28170 377922 28226
rect 377978 28170 408518 28226
rect 408574 28170 408642 28226
rect 408698 28170 439238 28226
rect 439294 28170 439362 28226
rect 439418 28170 469958 28226
rect 470014 28170 470082 28226
rect 470138 28170 500678 28226
rect 500734 28170 500802 28226
rect 500858 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 39878 28102
rect 39934 28046 40002 28102
rect 40058 28046 70598 28102
rect 70654 28046 70722 28102
rect 70778 28046 101318 28102
rect 101374 28046 101442 28102
rect 101498 28046 132038 28102
rect 132094 28046 132162 28102
rect 132218 28046 162758 28102
rect 162814 28046 162882 28102
rect 162938 28046 193478 28102
rect 193534 28046 193602 28102
rect 193658 28046 224198 28102
rect 224254 28046 224322 28102
rect 224378 28046 254918 28102
rect 254974 28046 255042 28102
rect 255098 28046 285638 28102
rect 285694 28046 285762 28102
rect 285818 28046 316358 28102
rect 316414 28046 316482 28102
rect 316538 28046 347078 28102
rect 347134 28046 347202 28102
rect 347258 28046 377798 28102
rect 377854 28046 377922 28102
rect 377978 28046 408518 28102
rect 408574 28046 408642 28102
rect 408698 28046 439238 28102
rect 439294 28046 439362 28102
rect 439418 28046 469958 28102
rect 470014 28046 470082 28102
rect 470138 28046 500678 28102
rect 500734 28046 500802 28102
rect 500858 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 39878 27978
rect 39934 27922 40002 27978
rect 40058 27922 70598 27978
rect 70654 27922 70722 27978
rect 70778 27922 101318 27978
rect 101374 27922 101442 27978
rect 101498 27922 132038 27978
rect 132094 27922 132162 27978
rect 132218 27922 162758 27978
rect 162814 27922 162882 27978
rect 162938 27922 193478 27978
rect 193534 27922 193602 27978
rect 193658 27922 224198 27978
rect 224254 27922 224322 27978
rect 224378 27922 254918 27978
rect 254974 27922 255042 27978
rect 255098 27922 285638 27978
rect 285694 27922 285762 27978
rect 285818 27922 316358 27978
rect 316414 27922 316482 27978
rect 316538 27922 347078 27978
rect 347134 27922 347202 27978
rect 347258 27922 377798 27978
rect 377854 27922 377922 27978
rect 377978 27922 408518 27978
rect 408574 27922 408642 27978
rect 408698 27922 439238 27978
rect 439294 27922 439362 27978
rect 439418 27922 469958 27978
rect 470014 27922 470082 27978
rect 470138 27922 500678 27978
rect 500734 27922 500802 27978
rect 500858 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use user_proj_example  mprj
timestamp 0
transform 1 0 20000 0 1 20000
box 914 0 499278 500000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 3154 -1644 3774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 21154 -1644 21774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 21154 520886 21774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 39154 -1644 39774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 39154 520886 39774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 57154 -1644 57774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 57154 520886 57774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 75154 -1644 75774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 75154 520886 75774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 93154 -1644 93774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 93154 520886 93774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 111154 -1644 111774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 111154 520886 111774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 -1644 129774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 520886 129774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 -1644 147774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 520886 147774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 -1644 165774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 520886 165774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 -1644 183774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 520886 183774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 -1644 201774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 520886 201774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 -1644 219774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 520886 219774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 -1644 237774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 520886 237774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 -1644 255774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 520886 255774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 -1644 273774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 520886 273774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 -1644 291774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 520886 291774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 -1644 309774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 520886 309774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 -1644 327774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 520886 327774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 -1644 345774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 520886 345774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 -1644 363774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 520886 363774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 -1644 381774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 520886 381774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 -1644 399774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 520886 399774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 -1644 417774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 520886 417774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 -1644 435774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 520886 435774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 -1644 453774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 520886 453774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 -1644 471774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 520886 471774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 -1644 489774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 520886 489774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 507154 -1644 507774 18186 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 507154 520886 507774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 525154 -1644 525774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 543154 -1644 543774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 561154 -1644 561774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 579154 -1644 579774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 6874 -1644 7494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 24874 -1644 25494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 24874 520886 25494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 42874 -1644 43494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 42874 520886 43494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 60874 -1644 61494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 60874 520886 61494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 78874 -1644 79494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 78874 520886 79494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96874 -1644 97494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96874 520886 97494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 -1644 115494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 520886 115494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 -1644 133494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 520886 133494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 -1644 151494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 520886 151494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 -1644 169494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 520886 169494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 -1644 187494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 520886 187494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 -1644 205494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 520886 205494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 -1644 223494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 520886 223494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 -1644 241494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 520886 241494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 -1644 259494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 520886 259494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 -1644 277494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 520886 277494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 -1644 295494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 520886 295494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 -1644 313494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 520886 313494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 -1644 331494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 520886 331494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 348874 -1644 349494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 348874 520886 349494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 -1644 367494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 520886 367494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 384874 -1644 385494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 384874 520886 385494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 -1644 403494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 520886 403494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 -1644 421494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 520886 421494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 -1644 439494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 520886 439494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 -1644 457494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 520886 457494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 474874 -1644 475494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 474874 520886 475494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 -1644 493494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 520886 493494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 510874 -1644 511494 18186 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 510874 520886 511494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 528874 -1644 529494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 546874 -1644 547494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 564874 -1644 565494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 582874 -1644 583494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 516190 508322 516190 508322 0 vdd
rlabel via4 500830 514322 500830 514322 0 vss
rlabel metal3 595098 7336 595098 7336 0 io_in[0]
rlabel metal3 594986 403816 594986 403816 0 io_in[10]
rlabel metal2 166978 519960 166978 519960 0 io_in[11]
rlabel metal3 594426 483112 594426 483112 0 io_in[12]
rlabel metal2 193942 519960 193942 519960 0 io_in[13]
rlabel metal3 595672 561624 595672 561624 0 io_in[14]
rlabel metal2 219870 519960 219870 519960 0 io_in[15]
rlabel metal2 233198 519960 233198 519960 0 io_in[16]
rlabel metal2 452312 593138 452312 593138 0 io_in[17]
rlabel metal2 259462 519960 259462 519960 0 io_in[18]
rlabel metal2 272510 519960 272510 519960 0 io_in[19]
rlabel metal3 594538 46984 594538 46984 0 io_in[1]
rlabel metal2 284914 519960 284914 519960 0 io_in[20]
rlabel metal3 188384 590184 188384 590184 0 io_in[21]
rlabel metal2 311178 519960 311178 519960 0 io_in[22]
rlabel metal2 54432 595672 54432 595672 0 io_in[23]
rlabel metal3 392 586712 392 586712 0 io_in[24]
rlabel metal3 392 544600 392 544600 0 io_in[25]
rlabel metal2 363594 519960 363594 519960 0 io_in[26]
rlabel metal3 392 459368 392 459368 0 io_in[27]
rlabel metal2 389970 519960 389970 519960 0 io_in[28]
rlabel metal3 392 375032 392 375032 0 io_in[29]
rlabel metal2 49798 519960 49798 519960 0 io_in[2]
rlabel metal3 4942 333368 4942 333368 0 io_in[30]
rlabel metal2 429114 519960 429114 519960 0 io_in[31]
rlabel metal2 442218 519960 442218 519960 0 io_in[32]
rlabel metal3 392 205520 392 205520 0 io_in[33]
rlabel metal3 392 163352 392 163352 0 io_in[34]
rlabel metal3 392 121184 392 121184 0 io_in[35]
rlabel metal2 494634 519960 494634 519960 0 io_in[36]
rlabel metal3 2310 36792 2310 36792 0 io_in[37]
rlabel metal3 594706 126280 594706 126280 0 io_in[3]
rlabel metal2 75726 519960 75726 519960 0 io_in[4]
rlabel metal3 594818 205576 594818 205576 0 io_in[5]
rlabel metal3 594874 245224 594874 245224 0 io_in[6]
rlabel metal2 115318 519960 115318 519960 0 io_in[7]
rlabel metal2 231896 525784 231896 525784 0 io_in[8]
rlabel metal2 141246 519960 141246 519960 0 io_in[9]
rlabel metal2 27258 519960 27258 519960 0 io_oeb[0]
rlabel metal2 523320 481544 523320 481544 0 io_oeb[10]
rlabel metal2 171570 519960 171570 519960 0 io_oeb[11]
rlabel metal2 184926 519960 184926 519960 0 io_oeb[12]
rlabel metal3 593250 548968 593250 548968 0 io_oeb[13]
rlabel metal2 211358 519960 211358 519960 0 io_oeb[14]
rlabel metal2 539896 595672 539896 595672 0 io_oeb[15]
rlabel metal2 237622 519960 237622 519960 0 io_oeb[16]
rlabel metal2 250446 519960 250446 519960 0 io_oeb[17]
rlabel metal2 263074 519960 263074 519960 0 io_oeb[18]
rlabel metal2 276178 519960 276178 519960 0 io_oeb[19]
rlabel metal3 594594 73416 594594 73416 0 io_oeb[1]
rlabel metal2 208936 595672 208936 595672 0 io_oeb[20]
rlabel metal2 143080 595672 143080 595672 0 io_oeb[21]
rlabel metal2 77336 572922 77336 572922 0 io_oeb[22]
rlabel metal2 328594 519960 328594 519960 0 io_oeb[23]
rlabel metal3 392 558320 392 558320 0 io_oeb[24]
rlabel metal3 2758 516824 2758 516824 0 io_oeb[25]
rlabel metal3 392 473984 392 473984 0 io_oeb[26]
rlabel metal2 381486 519960 381486 519960 0 io_oeb[27]
rlabel metal2 394114 519960 394114 519960 0 io_oeb[28]
rlabel metal2 407274 519960 407274 519960 0 io_oeb[29]
rlabel metal2 53886 519960 53886 519960 0 io_oeb[2]
rlabel metal3 1526 305144 1526 305144 0 io_oeb[30]
rlabel metal3 3262 262808 3262 262808 0 io_oeb[31]
rlabel metal2 447006 519960 447006 519960 0 io_oeb[32]
rlabel metal3 392 177128 392 177128 0 io_oeb[33]
rlabel metal2 472738 519960 472738 519960 0 io_oeb[34]
rlabel metal3 4830 93464 4830 93464 0 io_oeb[35]
rlabel metal3 1470 51128 1470 51128 0 io_oeb[36]
rlabel metal2 512806 519960 512806 519960 0 io_oeb[37]
rlabel metal2 538440 341096 538440 341096 0 io_oeb[3]
rlabel metal3 595672 191800 595672 191800 0 io_oeb[4]
rlabel metal2 541800 375648 541800 375648 0 io_oeb[5]
rlabel metal3 595672 270928 595672 270928 0 io_oeb[6]
rlabel metal2 119406 519960 119406 519960 0 io_oeb[7]
rlabel metal3 595672 350056 595672 350056 0 io_oeb[8]
rlabel metal2 145138 519960 145138 519960 0 io_oeb[9]
rlabel metal3 594482 20552 594482 20552 0 io_out[0]
rlabel metal2 163366 519960 163366 519960 0 io_out[10]
rlabel metal2 567000 492408 567000 492408 0 io_out[11]
rlabel metal2 189518 519960 189518 519960 0 io_out[12]
rlabel metal3 595672 534968 595672 534968 0 io_out[13]
rlabel metal2 215250 519960 215250 519960 0 io_out[14]
rlabel metal2 562632 593082 562632 593082 0 io_out[15]
rlabel metal2 241766 519960 241766 519960 0 io_out[16]
rlabel metal2 430136 568260 430136 568260 0 io_out[17]
rlabel metal2 335160 577976 335160 577976 0 io_out[18]
rlabel metal2 280770 519960 280770 519960 0 io_out[19]
rlabel metal2 44674 519960 44674 519960 0 io_out[1]
rlabel metal2 230888 595672 230888 595672 0 io_out[20]
rlabel metal3 166432 590184 166432 590184 0 io_out[21]
rlabel metal2 99176 571620 99176 571620 0 io_out[22]
rlabel metal2 333018 519960 333018 519960 0 io_out[23]
rlabel metal2 346290 519960 346290 519960 0 io_out[24]
rlabel metal2 359646 519960 359646 519960 0 io_out[25]
rlabel metal3 392 487760 392 487760 0 io_out[26]
rlabel metal3 392 445592 392 445592 0 io_out[27]
rlabel metal3 1582 403928 1582 403928 0 io_out[28]
rlabel metal2 411810 519960 411810 519960 0 io_out[29]
rlabel metal3 595672 99344 595672 99344 0 io_out[2]
rlabel metal2 425166 519960 425166 519960 0 io_out[30]
rlabel metal2 437794 519960 437794 519960 0 io_out[31]
rlabel metal3 392 233912 392 233912 0 io_out[32]
rlabel metal3 3206 192248 3206 192248 0 io_out[33]
rlabel metal2 477330 519960 477330 519960 0 io_out[34]
rlabel metal2 490686 519960 490686 519960 0 io_out[35]
rlabel metal3 392 64400 392 64400 0 io_out[36]
rlabel metal3 2702 22680 2702 22680 0 io_out[37]
rlabel metal2 70938 519960 70938 519960 0 io_out[3]
rlabel metal2 570360 364672 570360 364672 0 io_out[4]
rlabel metal2 97566 519960 97566 519960 0 io_out[5]
rlabel metal3 595672 257600 595672 257600 0 io_out[6]
rlabel metal2 123298 519960 123298 519960 0 io_out[7]
rlabel metal3 595672 336728 595672 336728 0 io_out[8]
rlabel metal3 595672 376712 595672 376712 0 io_out[9]
rlabel metal2 213192 3150 213192 3150 0 la_data_in[0]
rlabel metal2 270312 3990 270312 3990 0 la_data_in[10]
rlabel metal2 252728 14658 252728 14658 0 la_data_in[11]
rlabel metal2 281736 4102 281736 4102 0 la_data_in[12]
rlabel metal2 262136 18018 262136 18018 0 la_data_in[13]
rlabel metal2 266126 20104 266126 20104 0 la_data_in[14]
rlabel metal2 298088 392 298088 392 0 la_data_in[15]
rlabel metal2 304584 4158 304584 4158 0 la_data_in[16]
rlabel metal2 307608 6048 307608 6048 0 la_data_in[17]
rlabel metal2 288792 16408 288792 16408 0 la_data_in[18]
rlabel metal2 290360 18914 290360 18914 0 la_data_in[19]
rlabel metal2 218904 5726 218904 5726 0 la_data_in[1]
rlabel metal2 327432 4102 327432 4102 0 la_data_in[20]
rlabel metal2 333144 5670 333144 5670 0 la_data_in[21]
rlabel metal2 304262 20104 304262 20104 0 la_data_in[22]
rlabel metal2 309176 18858 309176 18858 0 la_data_in[23]
rlabel metal2 349832 392 349832 392 0 la_data_in[24]
rlabel metal2 355992 3262 355992 3262 0 la_data_in[25]
rlabel metal2 361704 3990 361704 3990 0 la_data_in[26]
rlabel metal2 327782 20104 327782 20104 0 la_data_in[27]
rlabel metal2 335384 15568 335384 15568 0 la_data_in[28]
rlabel metal2 378392 392 378392 392 0 la_data_in[29]
rlabel metal2 210392 15722 210392 15722 0 la_data_in[2]
rlabel metal2 384552 4102 384552 4102 0 la_data_in[30]
rlabel metal2 374136 16128 374136 16128 0 la_data_in[31]
rlabel metal3 355936 16856 355936 16856 0 la_data_in[32]
rlabel metal2 401688 3262 401688 3262 0 la_data_in[33]
rlabel metal2 360920 15554 360920 15554 0 la_data_in[34]
rlabel metal2 365624 14770 365624 14770 0 la_data_in[35]
rlabel metal2 418824 3206 418824 3206 0 la_data_in[36]
rlabel metal2 375704 15512 375704 15512 0 la_data_in[37]
rlabel metal2 383544 14952 383544 14952 0 la_data_in[38]
rlabel metal2 383726 20104 383726 20104 0 la_data_in[39]
rlabel metal2 215166 20104 215166 20104 0 la_data_in[3]
rlabel metal3 410004 7896 410004 7896 0 la_data_in[40]
rlabel metal2 447384 3374 447384 3374 0 la_data_in[41]
rlabel metal2 398552 18914 398552 18914 0 la_data_in[42]
rlabel metal2 403256 19026 403256 19026 0 la_data_in[43]
rlabel metal2 407960 19138 407960 19138 0 la_data_in[44]
rlabel metal2 470232 5894 470232 5894 0 la_data_in[45]
rlabel metal2 475664 392 475664 392 0 la_data_in[46]
rlabel metal2 422072 17402 422072 17402 0 la_data_in[47]
rlabel metal2 426776 18970 426776 18970 0 la_data_in[48]
rlabel metal2 493080 3262 493080 3262 0 la_data_in[49]
rlabel metal2 235592 392 235592 392 0 la_data_in[4]
rlabel metal2 498792 4214 498792 4214 0 la_data_in[50]
rlabel metal2 504224 392 504224 392 0 la_data_in[51]
rlabel metal2 445438 20104 445438 20104 0 la_data_in[52]
rlabel metal2 515928 3318 515928 3318 0 la_data_in[53]
rlabel metal2 521192 392 521192 392 0 la_data_in[54]
rlabel metal2 526568 392 526568 392 0 la_data_in[55]
rlabel metal2 533064 3262 533064 3262 0 la_data_in[56]
rlabel metal2 538160 392 538160 392 0 la_data_in[57]
rlabel metal2 473816 18466 473816 18466 0 la_data_in[58]
rlabel metal2 478520 17234 478520 17234 0 la_data_in[59]
rlabel metal2 240968 392 240968 392 0 la_data_in[5]
rlabel metal2 555128 392 555128 392 0 la_data_in[60]
rlabel metal2 561176 2688 561176 2688 0 la_data_in[61]
rlabel metal2 567336 3990 567336 3990 0 la_data_in[62]
rlabel metal2 497336 18018 497336 18018 0 la_data_in[63]
rlabel metal2 247184 392 247184 392 0 la_data_in[6]
rlabel metal2 233912 17458 233912 17458 0 la_data_in[7]
rlabel metal3 258384 4200 258384 4200 0 la_data_in[8]
rlabel metal2 264600 3262 264600 3262 0 la_data_in[9]
rlabel metal2 215096 5670 215096 5670 0 la_data_out[0]
rlabel metal2 272216 2366 272216 2366 0 la_data_out[10]
rlabel metal2 277928 3206 277928 3206 0 la_data_out[11]
rlabel metal3 262752 3976 262752 3976 0 la_data_out[12]
rlabel metal2 289352 3150 289352 3150 0 la_data_out[13]
rlabel metal2 295064 2534 295064 2534 0 la_data_out[14]
rlabel metal2 275464 15792 275464 15792 0 la_data_out[15]
rlabel metal2 306096 392 306096 392 0 la_data_out[16]
rlabel metal2 312200 2646 312200 2646 0 la_data_out[17]
rlabel metal2 286454 20104 286454 20104 0 la_data_out[18]
rlabel metal2 306936 15288 306936 15288 0 la_data_out[19]
rlabel metal2 207256 15834 207256 15834 0 la_data_out[1]
rlabel metal2 329336 7350 329336 7350 0 la_data_out[20]
rlabel metal2 334656 392 334656 392 0 la_data_out[21]
rlabel metal2 306040 14658 306040 14658 0 la_data_out[22]
rlabel metal2 312424 13944 312424 13944 0 la_data_out[23]
rlabel metal2 351624 392 351624 392 0 la_data_out[24]
rlabel metal2 357896 4886 357896 4886 0 la_data_out[25]
rlabel metal2 363608 1470 363608 1470 0 la_data_out[26]
rlabel metal2 329560 18018 329560 18018 0 la_data_out[27]
rlabel metal2 334264 15498 334264 15498 0 la_data_out[28]
rlabel metal2 380744 4158 380744 4158 0 la_data_out[29]
rlabel metal2 211960 15778 211960 15778 0 la_data_out[2]
rlabel metal2 352744 15848 352744 15848 0 la_data_out[30]
rlabel metal2 349496 16464 349496 16464 0 la_data_out[31]
rlabel metal2 397152 392 397152 392 0 la_data_out[32]
rlabel metal2 357784 14658 357784 14658 0 la_data_out[33]
rlabel metal2 408744 392 408744 392 0 la_data_out[34]
rlabel metal2 367976 17024 367976 17024 0 la_data_out[35]
rlabel metal2 420728 1526 420728 1526 0 la_data_out[36]
rlabel metal2 425768 392 425768 392 0 la_data_out[37]
rlabel metal2 379736 8036 379736 8036 0 la_data_out[38]
rlabel metal2 407624 14560 407624 14560 0 la_data_out[39]
rlabel metal2 232008 392 232008 392 0 la_data_out[3]
rlabel metal2 443576 7462 443576 7462 0 la_data_out[40]
rlabel metal2 449288 4886 449288 4886 0 la_data_out[41]
rlabel metal2 454272 392 454272 392 0 la_data_out[42]
rlabel metal2 404824 17234 404824 17234 0 la_data_out[43]
rlabel metal2 465864 392 465864 392 0 la_data_out[44]
rlabel metal2 472136 3150 472136 3150 0 la_data_out[45]
rlabel metal2 477848 5838 477848 5838 0 la_data_out[46]
rlabel metal2 423640 16338 423640 16338 0 la_data_out[47]
rlabel metal2 426776 5516 426776 5516 0 la_data_out[48]
rlabel metal2 494984 5670 494984 5670 0 la_data_out[49]
rlabel metal2 237384 392 237384 392 0 la_data_out[4]
rlabel metal2 500696 3990 500696 3990 0 la_data_out[50]
rlabel metal2 506408 1470 506408 1470 0 la_data_out[51]
rlabel metal2 447006 20104 447006 20104 0 la_data_out[52]
rlabel metal2 517608 392 517608 392 0 la_data_out[53]
rlabel metal2 522984 392 522984 392 0 la_data_out[54]
rlabel metal2 529256 5726 529256 5726 0 la_data_out[55]
rlabel metal2 465976 15610 465976 15610 0 la_data_out[56]
rlabel metal2 539952 392 539952 392 0 la_data_out[57]
rlabel metal2 546392 1582 546392 1582 0 la_data_out[58]
rlabel metal2 480088 14658 480088 14658 0 la_data_out[59]
rlabel metal2 226072 17178 226072 17178 0 la_data_out[5]
rlabel metal2 484792 16338 484792 16338 0 la_data_out[60]
rlabel metal2 563136 392 563136 392 0 la_data_out[61]
rlabel metal2 494200 15442 494200 15442 0 la_data_out[62]
rlabel metal2 498904 19138 498904 19138 0 la_data_out[63]
rlabel metal2 249032 392 249032 392 0 la_data_out[6]
rlabel metal2 235480 17514 235480 17514 0 la_data_out[7]
rlabel metal2 260792 2422 260792 2422 0 la_data_out[8]
rlabel metal2 266504 2254 266504 2254 0 la_data_out[9]
rlabel metal2 217000 5838 217000 5838 0 la_oenb[0]
rlabel metal2 274120 2590 274120 2590 0 la_oenb[10]
rlabel metal2 279832 2198 279832 2198 0 la_oenb[11]
rlabel metal2 260568 18858 260568 18858 0 la_oenb[12]
rlabel metal2 264502 20104 264502 20104 0 la_oenb[13]
rlabel metal2 296968 2310 296968 2310 0 la_oenb[14]
rlabel metal2 302680 2422 302680 2422 0 la_oenb[15]
rlabel metal2 308392 2702 308392 2702 0 la_oenb[16]
rlabel metal2 283990 20104 283990 20104 0 la_oenb[17]
rlabel metal2 288792 18858 288792 18858 0 la_oenb[18]
rlabel metal2 325528 3150 325528 3150 0 la_oenb[19]
rlabel metal2 208824 15610 208824 15610 0 la_oenb[1]
rlabel metal2 331240 2590 331240 2590 0 la_oenb[20]
rlabel metal2 336952 2310 336952 2310 0 la_oenb[21]
rlabel metal2 307510 20104 307510 20104 0 la_oenb[22]
rlabel metal2 311542 20104 311542 20104 0 la_oenb[23]
rlabel metal2 354088 3150 354088 3150 0 la_oenb[24]
rlabel metal2 359800 2422 359800 2422 0 la_oenb[25]
rlabel metal2 326424 18970 326424 18970 0 la_oenb[26]
rlabel metal2 331030 20104 331030 20104 0 la_oenb[27]
rlabel metal2 376936 3318 376936 3318 0 la_oenb[28]
rlabel metal2 382648 2310 382648 2310 0 la_oenb[29]
rlabel metal2 213430 20104 213430 20104 0 la_oenb[2]
rlabel metal2 388248 4200 388248 4200 0 la_oenb[30]
rlabel metal2 349944 15610 349944 15610 0 la_oenb[31]
rlabel metal2 399896 3150 399896 3150 0 la_oenb[32]
rlabel metal2 405160 392 405160 392 0 la_oenb[33]
rlabel metal2 411208 1694 411208 1694 0 la_oenb[34]
rlabel metal3 415520 5432 415520 5432 0 la_oenb[35]
rlabel metal2 422128 392 422128 392 0 la_oenb[36]
rlabel metal2 378168 17178 378168 17178 0 la_oenb[37]
rlabel metal2 382872 19026 382872 19026 0 la_oenb[38]
rlabel metal2 439768 1470 439768 1470 0 la_oenb[39]
rlabel metal2 233800 392 233800 392 0 la_oenb[3]
rlabel metal2 445368 4200 445368 4200 0 la_oenb[40]
rlabel metal2 450688 392 450688 392 0 la_oenb[41]
rlabel metal2 401688 18858 401688 18858 0 la_oenb[42]
rlabel metal2 406392 14658 406392 14658 0 la_oenb[43]
rlabel metal2 468328 1582 468328 1582 0 la_oenb[44]
rlabel metal2 474040 3318 474040 3318 0 la_oenb[45]
rlabel metal2 427336 14896 427336 14896 0 la_oenb[46]
rlabel metal2 425264 56 425264 56 0 la_oenb[47]
rlabel metal2 490896 392 490896 392 0 la_oenb[48]
rlabel metal3 491400 7840 491400 7840 0 la_oenb[49]
rlabel metal2 239176 392 239176 392 0 la_oenb[4]
rlabel metal2 439320 19138 439320 19138 0 la_oenb[50]
rlabel metal2 444024 19082 444024 19082 0 la_oenb[51]
rlabel metal2 448728 19026 448728 19026 0 la_oenb[52]
rlabel metal2 519736 1638 519736 1638 0 la_oenb[53]
rlabel metal2 525448 4158 525448 4158 0 la_oenb[54]
rlabel metal2 531160 2590 531160 2590 0 la_oenb[55]
rlabel metal2 467278 20104 467278 20104 0 la_oenb[56]
rlabel metal2 542696 2534 542696 2534 0 la_oenb[57]
rlabel metal2 548296 2478 548296 2478 0 la_oenb[58]
rlabel metal2 496440 12824 496440 12824 0 la_oenb[59]
rlabel metal2 227640 17290 227640 17290 0 la_oenb[5]
rlabel metal2 559720 2422 559720 2422 0 la_oenb[60]
rlabel metal2 565432 2366 565432 2366 0 la_oenb[61]
rlabel metal2 495768 19082 495768 19082 0 la_oenb[62]
rlabel metal2 499702 20104 499702 20104 0 la_oenb[63]
rlabel metal2 232344 17402 232344 17402 0 la_oenb[6]
rlabel metal2 257096 2534 257096 2534 0 la_oenb[7]
rlabel metal2 262696 2478 262696 2478 0 la_oenb[8]
rlabel metal2 267736 392 267736 392 0 la_oenb[9]
rlabel metal2 502040 18970 502040 18970 0 user_irq[0]
rlabel metal2 581896 392 581896 392 0 user_irq[1]
rlabel metal3 580776 4760 580776 4760 0 user_irq[2]
rlabel metal2 11592 3990 11592 3990 0 wb_clk_i
rlabel metal2 13384 5670 13384 5670 0 wb_rst_i
rlabel metal2 15176 6510 15176 6510 0 wbs_ack_o
rlabel metal2 23016 3150 23016 3150 0 wbs_adr_i[0]
rlabel metal2 97496 18858 97496 18858 0 wbs_adr_i[10]
rlabel metal2 92792 392 92792 392 0 wbs_adr_i[11]
rlabel metal2 98280 392 98280 392 0 wbs_adr_i[12]
rlabel metal2 104384 392 104384 392 0 wbs_adr_i[13]
rlabel metal2 116102 20104 116102 20104 0 wbs_adr_i[14]
rlabel metal2 121016 18522 121016 18522 0 wbs_adr_i[15]
rlabel metal2 121352 392 121352 392 0 wbs_adr_i[16]
rlabel metal2 126728 392 126728 392 0 wbs_adr_i[17]
rlabel metal2 132944 392 132944 392 0 wbs_adr_i[18]
rlabel metal2 138376 392 138376 392 0 wbs_adr_i[19]
rlabel metal2 30408 8190 30408 8190 0 wbs_adr_i[1]
rlabel metal2 144606 20104 144606 20104 0 wbs_adr_i[20]
rlabel metal2 148526 20104 148526 20104 0 wbs_adr_i[21]
rlabel metal3 154504 4312 154504 4312 0 wbs_adr_i[22]
rlabel metal2 161784 2590 161784 2590 0 wbs_adr_i[23]
rlabel metal3 165256 4312 165256 4312 0 wbs_adr_i[24]
rlabel metal2 168056 12418 168056 12418 0 wbs_adr_i[25]
rlabel metal2 172046 20104 172046 20104 0 wbs_adr_i[26]
rlabel metal3 180544 6440 180544 6440 0 wbs_adr_i[27]
rlabel metal2 190344 3262 190344 3262 0 wbs_adr_i[28]
rlabel metal3 191296 6328 191296 6328 0 wbs_adr_i[29]
rlabel metal2 37464 392 37464 392 0 wbs_adr_i[2]
rlabel metal2 191576 12194 191576 12194 0 wbs_adr_i[30]
rlabel metal2 195566 20104 195566 20104 0 wbs_adr_i[31]
rlabel metal2 45864 6006 45864 6006 0 wbs_adr_i[3]
rlabel metal2 53480 5670 53480 5670 0 wbs_adr_i[4]
rlabel metal2 74158 20104 74158 20104 0 wbs_adr_i[5]
rlabel metal2 78302 20104 78302 20104 0 wbs_adr_i[6]
rlabel metal2 69608 392 69608 392 0 wbs_adr_i[7]
rlabel metal2 75824 392 75824 392 0 wbs_adr_i[8]
rlabel metal2 92582 20104 92582 20104 0 wbs_adr_i[9]
rlabel metal2 17304 2310 17304 2310 0 wbs_cyc_i
rlabel metal2 24920 2478 24920 2478 0 wbs_dat_i[0]
rlabel metal2 98686 20104 98686 20104 0 wbs_dat_i[10]
rlabel metal2 94584 392 94584 392 0 wbs_dat_i[11]
rlabel metal2 100856 9030 100856 9030 0 wbs_dat_i[12]
rlabel metal2 106176 392 106176 392 0 wbs_dat_i[13]
rlabel metal2 117726 20104 117726 20104 0 wbs_dat_i[14]
rlabel metal2 117768 392 117768 392 0 wbs_dat_i[15]
rlabel metal2 123200 392 123200 392 0 wbs_dat_i[16]
rlabel metal2 131670 20104 131670 20104 0 wbs_dat_i[17]
rlabel metal2 134792 392 134792 392 0 wbs_dat_i[18]
rlabel metal2 140112 392 140112 392 0 wbs_dat_i[19]
rlabel metal2 51646 20104 51646 20104 0 wbs_dat_i[1]
rlabel metal3 145656 4648 145656 4648 0 wbs_dat_i[20]
rlabel metal3 150920 4312 150920 4312 0 wbs_dat_i[21]
rlabel metal3 156296 4648 156296 4648 0 wbs_dat_i[22]
rlabel metal2 163688 2646 163688 2646 0 wbs_dat_i[23]
rlabel metal3 167048 4088 167048 4088 0 wbs_dat_i[24]
rlabel metal2 168854 20104 168854 20104 0 wbs_dat_i[25]
rlabel metal3 176960 5096 176960 5096 0 wbs_dat_i[26]
rlabel metal2 186536 3094 186536 3094 0 wbs_dat_i[27]
rlabel metal2 192248 3318 192248 3318 0 wbs_dat_i[28]
rlabel metal3 188440 5992 188440 5992 0 wbs_dat_i[29]
rlabel metal2 39256 392 39256 392 0 wbs_dat_i[2]
rlabel metal2 192374 20104 192374 20104 0 wbs_dat_i[30]
rlabel metal2 209384 3374 209384 3374 0 wbs_dat_i[31]
rlabel metal2 47768 5838 47768 5838 0 wbs_dat_i[3]
rlabel metal2 55384 5894 55384 5894 0 wbs_dat_i[4]
rlabel metal2 75166 20104 75166 20104 0 wbs_dat_i[5]
rlabel metal2 66024 392 66024 392 0 wbs_dat_i[6]
rlabel metal2 72408 6846 72408 6846 0 wbs_dat_i[7]
rlabel metal2 77616 392 77616 392 0 wbs_dat_i[8]
rlabel metal2 94262 20104 94262 20104 0 wbs_dat_i[9]
rlabel metal2 26824 2422 26824 2422 0 wbs_dat_o[0]
rlabel metal2 91000 392 91000 392 0 wbs_dat_o[10]
rlabel metal2 96432 392 96432 392 0 wbs_dat_o[11]
rlabel metal2 109662 20104 109662 20104 0 wbs_dat_o[12]
rlabel metal2 114590 20104 114590 20104 0 wbs_dat_o[13]
rlabel metal2 119350 20104 119350 20104 0 wbs_dat_o[14]
rlabel metal2 119560 392 119560 392 0 wbs_dat_o[15]
rlabel metal2 124936 392 124936 392 0 wbs_dat_o[16]
rlabel metal2 133182 20104 133182 20104 0 wbs_dat_o[17]
rlabel metal2 138110 20104 138110 20104 0 wbs_dat_o[18]
rlabel metal2 142870 20104 142870 20104 0 wbs_dat_o[19]
rlabel metal2 53214 20104 53214 20104 0 wbs_dat_o[1]
rlabel metal3 147336 4312 147336 4312 0 wbs_dat_o[20]
rlabel metal3 152712 4200 152712 4200 0 wbs_dat_o[21]
rlabel metal3 158088 4200 158088 4200 0 wbs_dat_o[22]
rlabel metal3 163464 4200 163464 4200 0 wbs_dat_o[23]
rlabel metal3 168896 4536 168896 4536 0 wbs_dat_o[24]
rlabel metal2 170422 20104 170422 20104 0 wbs_dat_o[25]
rlabel metal3 178752 6216 178752 6216 0 wbs_dat_o[26]
rlabel metal2 188440 3150 188440 3150 0 wbs_dat_o[27]
rlabel metal3 189504 5096 189504 5096 0 wbs_dat_o[28]
rlabel metal2 189910 20104 189910 20104 0 wbs_dat_o[29]
rlabel metal2 41104 392 41104 392 0 wbs_dat_o[2]
rlabel metal2 193942 20104 193942 20104 0 wbs_dat_o[30]
rlabel metal2 211288 3262 211288 3262 0 wbs_dat_o[31]
rlabel metal2 49672 5950 49672 5950 0 wbs_dat_o[3]
rlabel metal2 72310 20104 72310 20104 0 wbs_dat_o[4]
rlabel metal2 76734 20104 76734 20104 0 wbs_dat_o[5]
rlabel metal2 67816 392 67816 392 0 wbs_dat_o[6]
rlabel metal2 74200 6790 74200 6790 0 wbs_dat_o[7]
rlabel metal2 91070 20104 91070 20104 0 wbs_dat_o[8]
rlabel metal2 95830 20104 95830 20104 0 wbs_dat_o[9]
rlabel metal2 28728 2534 28728 2534 0 wbs_sel_i[0]
rlabel metal2 54782 20104 54782 20104 0 wbs_sel_i[1]
rlabel metal2 43960 5726 43960 5726 0 wbs_sel_i[2]
rlabel metal2 51576 5782 51576 5782 0 wbs_sel_i[3]
rlabel metal2 18704 392 18704 392 0 wbs_stb_i
rlabel metal2 21112 2366 21112 2366 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
