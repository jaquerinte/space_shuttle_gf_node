// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
//-----------------------------------------------------
// Project Name : a.out
// Function     : Main processor 
// Description  : This is the main processor
// Coder        : Jaquer AND VORIXO

//***Headers***
//***Module***
module parity_calculator #(
        parameter integer WORD_SIZE = 32,
        parameter integer ECCBITS = 7
    )
    (
        `ifdef USE_POWER_PINS
        inout wire vdda1,	// User area 1 3.3V supply
        inout wire vdda2,	// User area 2 3.3V supply
        inout wire vssa1,	// User area 1 analog ground
        inout wire vssa2,	// User area 2 analog ground
        inout wire vccd1,	// User area 1 1.8V supply
        inout wire vccd2,	// User area 2 1.8v supply
        inout wire vssd1,	// User area 1 digital ground
        inout wire vssd2,	// User area 2 digital ground
        `endif
        input  wire [WORD_SIZE - 1 : 0] data_to_register_i ,
        input  wire operate_i ,
        input  wire [2 : 0] operation_type_i,
        output wire [WORD_SIZE  + ECCBITS- 1 : 0] data_to_register_o 
    );

//***Internal logic generated by compiler***  
    wire intermidate_partity_bits [ECCBITS - 2 : 0];
    reg last_bit_value;
    reg intermidate_partity_bits_last;

//***Dumped Internal logic***
    assign  intermidate_partity_bits[0] = operate_i ?  data_to_register_i[0] ^ data_to_register_i[1] ^ data_to_register_i[3] ^ data_to_register_i[4]^ data_to_register_i[6]^ data_to_register_i[8]^ data_to_register_i[10]^ data_to_register_i[11]^ data_to_register_i[13]^ data_to_register_i[15]^ data_to_register_i[17]^ data_to_register_i[19]^ data_to_register_i[21]^ data_to_register_i[23] ^ data_to_register_i[25] ^ data_to_register_i[26]^ data_to_register_i[28]^ data_to_register_i[30] : 1'b0;
    assign  intermidate_partity_bits[1] = operate_i ?  data_to_register_i[0] ^ data_to_register_i[2] ^ data_to_register_i[3] ^ data_to_register_i[5]^ data_to_register_i[6]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[12]^ data_to_register_i[13]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[24] ^ data_to_register_i[25] ^ data_to_register_i[27]^ data_to_register_i[28]^ data_to_register_i[31] : 1'b0;
    assign  intermidate_partity_bits[2] = operate_i ?  data_to_register_i[1] ^ data_to_register_i[2] ^ data_to_register_i[3] ^ data_to_register_i[7]^ data_to_register_i[8]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[14]^ data_to_register_i[15]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24] ^ data_to_register_i[25] ^ data_to_register_i[29]^ data_to_register_i[30]^ data_to_register_i[31] : 1'b0;
    assign  intermidate_partity_bits[3] = operate_i ?  data_to_register_i[4] ^ data_to_register_i[5] ^ data_to_register_i[6] ^ data_to_register_i[7]^ data_to_register_i[8]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[18]^ data_to_register_i[19]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24] ^ data_to_register_i[25] : 1'b0;
    assign  intermidate_partity_bits[4] = operate_i ?  data_to_register_i[11] ^ data_to_register_i[12] ^ data_to_register_i[13] ^ data_to_register_i[14]^ data_to_register_i[15]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[18]^ data_to_register_i[19]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24]^ data_to_register_i[25]: 1'b0;
    assign  intermidate_partity_bits[5] = operate_i ?  data_to_register_i[26] ^ data_to_register_i[27] ^ data_to_register_i[28] ^ data_to_register_i[29]^ data_to_register_i[30]^ data_to_register_i[31]: 1'b0;
    //assign  intermidate_partity_bits[6] = operate_i ?  data_to_register_i[0] ^ data_to_register_i[1] ^ data_to_register_i[2] ^ data_to_register_i[3] ^ data_to_register_i[4]^ data_to_register_i[5]^ data_to_register_i[6]^ data_to_register_i[7]^ data_to_register_i[8]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[11]^ data_to_register_i[12]^ data_to_register_i[13]^ data_to_register_i[14]^ data_to_register_i[15]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[18]^ data_to_register_i[19]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24]^ data_to_register_i[25]^ data_to_register_i[26]^ data_to_register_i[27]^ data_to_register_i[28]^ data_to_register_i[29]^ data_to_register_i[30]^ data_to_register_i[31]: 1'b0;
    
    always @(*) begin
        intermidate_partity_bits_last = operate_i ?  data_to_register_i[0] ^ data_to_register_i[1] ^ data_to_register_i[2] ^ data_to_register_i[3] ^ data_to_register_i[4]^ data_to_register_i[5]^ data_to_register_i[6]^ data_to_register_i[7]^ data_to_register_i[8]^ data_to_register_i[9]^ data_to_register_i[10]^ data_to_register_i[11]^ data_to_register_i[12]^ data_to_register_i[13]^ data_to_register_i[14]^ data_to_register_i[15]^ data_to_register_i[16]^ data_to_register_i[17]^ data_to_register_i[18]^ data_to_register_i[19]^ data_to_register_i[20]^ data_to_register_i[21]^ data_to_register_i[22]^ data_to_register_i[23]^ data_to_register_i[24]^ data_to_register_i[25]^ data_to_register_i[26]^ data_to_register_i[27]^ data_to_register_i[28]^ data_to_register_i[29]^ data_to_register_i[30]^ data_to_register_i[31]: 1'b0;
        last_bit_value = intermidate_partity_bits_last ^ intermidate_partity_bits[0] ^ intermidate_partity_bits[1] ^ intermidate_partity_bits[2] ^ intermidate_partity_bits[3] ^ intermidate_partity_bits[4] ^ intermidate_partity_bits[5]  ; 
    end
    assign data_to_register_o = operation_type_i[2] == 1'b1 ?  {7'b0 ,data_to_register_i} : operation_type_i[0] == 1'b1 ? {7'b0 ,data_to_register_i}:{last_bit_value,data_to_register_i[31],data_to_register_i[30],data_to_register_i[29],data_to_register_i[28],data_to_register_i[27],data_to_register_i[26],intermidate_partity_bits[5],data_to_register_i[25],data_to_register_i[24],data_to_register_i[23],data_to_register_i[22],data_to_register_i[21],data_to_register_i[20],data_to_register_i[19],data_to_register_i[18],data_to_register_i[17],data_to_register_i[16],data_to_register_i[15],data_to_register_i[14],data_to_register_i[13],data_to_register_i[12],data_to_register_i[11],intermidate_partity_bits[4],data_to_register_i[10],data_to_register_i[9],data_to_register_i[8],data_to_register_i[7],data_to_register_i[6],data_to_register_i[5],data_to_register_i[4],intermidate_partity_bits[3],data_to_register_i[3],data_to_register_i[2],data_to_register_i[1],intermidate_partity_bits[2],data_to_register_i[0], intermidate_partity_bits[1], intermidate_partity_bits[0]};
    
//***Handcrafted Internal logic*** 
//TODO
endmodule
